* SPICE3 file created from amp-cs.ext - technology: sky130A

X0 A A A w_n15748_5772# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.791e+07u l=1e+06u
X1 A A A w_n15748_5772# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.791e+07u l=1e+06u
X2 A A A w_n15748_5772# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.791e+07u l=1e+06u
X3 A A A w_n15748_5772# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.791e+07u l=1e+06u
X4 A A A w_n15748_5772# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.791e+07u l=1e+06u
X5 A A A w_n15748_5772# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.791e+07u l=1e+06u
X6 A IN A VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8.6e+06u l=1e+06u
X7 A A A w_n15748_5772# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.79e+07u l=1e+06u
X8 A IN A VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8.6e+06u l=1e+06u
X9 A A A w_n15748_5772# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.791e+07u l=1e+06u
X10 A A A w_n15748_5772# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.79e+07u l=1e+06u
X11 A A A w_n15748_5772# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.791e+07u l=1e+06u
X12 A A A w_n15748_5772# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.791e+07u l=1e+06u
X13 A IN A VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8.6e+06u l=1e+06u
X14 A A A w_n15748_5772# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.791e+07u l=1e+06u
X15 A A A w_n15748_5772# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.791e+07u l=1e+06u
X16 A A A w_n15748_5772# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.791e+07u l=1e+06u
X17 A A A w_n15748_5772# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.791e+07u l=1e+06u
X18 A IN A VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8.6e+06u l=1e+06u
X19 A A A w_n15748_5772# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.791e+07u l=1e+06u
X20 A A A w_n15748_5772# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.791e+07u l=1e+06u
X21 A IN A VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8.6e+06u l=1e+06u
X22 A A A w_n15748_5772# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.791e+07u l=1e+06u
X23 A A A w_n15748_5772# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.791e+07u l=1e+06u
X24 A A A w_n15748_5772# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.791e+07u l=1e+06u
C0 A IN 1.92fF
C1 IN w_n15748_5772# 11.75fF
C2 A w_n15748_5772# 133.60fF
