*AMPLIFIER COMMON SOURCE


.subckt	ampcs_post	IN	OUT	Vd	GND
*label drain   gate    source  bulk    model           width   length
M1	OUT	IN	GND	GND	nshort_model	W=43u	L=1u
M2      OUT	A	Vd	Vd	pshort_model	W=479u  L=1u
M3      A	A	Vd	Vd	pshort_model	W=479u	L=1u

*parastics
R0 A.n14 A.t27 1513.26
R1 A.n5 A.t2 1509.02
R2 A.n22 A.t23 1296.1
R3 A.n14 A.t29 1295.86
R4 A.n15 A.t24 1295.86
R5 A.n16 A.t20 1295.86
R6 A.n17 A.t26 1295.86
R7 A.n18 A.t25 1295.86
R8 A.n19 A.t21 1295.86
R9 A.n20 A.t22 1295.86
R10 A.n21 A.t28 1295.86
R11 A.n13 A.t8 1294.89
R12 A.n12 A.t10 1294.89
R13 A.n11 A.t6 1294.89
R14 A.n10 A.t4 1294.89
R15 A.n9 A.t12 1294.89
R16 A.n8 A.t16 1294.89
R17 A.n7 A.t14 1294.89
R18 A.n6 A.t0 1294.89
R19 A.n5 A.t18 1294.43
R20 A.n44 A.t3 485.682
R21 A.n23 A.n13 467.459
R22 A.n23 A.n22 362.204
R23 A.n15 A.n14 214.49
R24 A.n16 A.n15 214.49
R25 A.n17 A.n16 214.49
R26 A.n18 A.n17 214.49
R27 A.n19 A.n18 214.49
R28 A.n20 A.n19 214.49
R29 A.n21 A.n20 214.49
R30 A.n22 A.n21 214.49
R31 A.n13 A.n12 210.284
R32 A.n12 A.n11 210.284
R33 A.n11 A.n10 210.284
R34 A.n10 A.n9 210.284
R35 A.n9 A.n8 210.284
R36 A.n8 A.n7 210.284
R37 A.n7 A.n6 210.284
R38 A.n6 A.n5 210.281
R39 A.n48 A.n47 108.702
R40 A.n47 A.n46 108.702
R41 A.n45 A.n44 108.458
R42 A.n46 A.n45 106.601
R43 A.n45 A.n3 102.663
R44 A.n46 A.n2 102.34
R45 A.n44 A.n4 102.339
R46 A.n47 A.n1 102.024
R47 A.n48 A.n0 101.714
R48 A A.n49 90.89
R49 A.n49 A.n48 88.446
R50 A.n25 A.n24 9.142
R51 A.n31 A.t7 8.161
R52 A.n35 A.t13 8.161
R53 A.n39 A.t15 8.161
R54 A.n43 A.t19 8.161
R55 A.n26 A.t9 7.915
R56 A.n28 A.t11 5.818
R57 A.n32 A.t5 5.818
R58 A.n36 A.t17 5.818
R59 A.n40 A.t1 5.818
R60 A.n0 A.n27 0.247
R61 A.n49 A.n23 0.196
R62 A.n27 A.n26 0.082
R63 A.n1 A.n31 0.082
R64 A.n2 A.n35 0.082
R65 A.n3 A.n39 0.082
R66 A.n4 A.n43 0.082
R67 A.n30 A.n29 0.044
R68 A.n34 A.n33 0.044
R69 A.n38 A.n37 0.044
R70 A.n42 A.n41 0.044
R71 A.n4 A.n42 0.042
R72 A.n3 A.n38 0.042
R73 A.n2 A.n34 0.042
R74 A.n1 A.n30 0.042
R75 A.n0 A.n25 0.042
R76 A.n29 A.n28 0.039
R77 A.n33 A.n32 0.039
R78 A.n37 A.n36 0.039
R79 A.n41 A.n40 0.039
R80 OUT.n13 OUT.t14 485.682
R81 OUT.n23 OUT.n2 210.416
R82 OUT.n32 OUT.t2 183.457
R83 OUT.n32 OUT.n30 160.642
R84 OUT.n28 OUT.n23 108.702
R85 OUT.n14 OUT.n13 108.458
R86 OUT.n14 OUT.n0 102.663
R87 OUT.n28 OUT.n4 102.34
R88 OUT.n13 OUT.n1 102.339
R89 OUT.n23 OUT.n3 102.024
R90 OUT.n32 OUT.n31 61.171
R91 OUT.n29 OUT.n14 56.73
R92 OUT OUT.n29 49.506
R93 OUT OUT.n32 49.353
R94 OUT.n29 OUT.n28 35.868
R95 OUT.n31 OUT.t4 26.093
R96 OUT.n31 OUT.t3 22.463
R97 OUT.n30 OUT.t1 21.625
R98 OUT.n30 OUT.t0 19.255
R99 OUT.n20 OUT.n19 9.142
R100 OUT.n8 OUT.t6 8.161
R101 OUT.n12 OUT.t10 8.161
R102 OUT.n18 OUT.t11 8.161
R103 OUT.n27 OUT.t9 8.161
R104 OUT.n21 OUT.t13 7.915
R105 OUT.n5 OUT.t12 5.818
R106 OUT.n9 OUT.t7 5.818
R107 OUT.n15 OUT.t8 5.818
R108 OUT.n24 OUT.t5 5.818
R109 OUT.n2 OUT.n22 0.247
R110 OUT.n22 OUT.n21 0.082
R111 OUT.n0 OUT.n8 0.082
R112 OUT.n1 OUT.n12 0.082
R113 OUT.n3 OUT.n18 0.082
R114 OUT.n4 OUT.n27 0.082
R115 OUT.n7 OUT.n6 0.044
R116 OUT.n11 OUT.n10 0.044
R117 OUT.n17 OUT.n16 0.044
R118 OUT.n26 OUT.n25 0.044
R119 OUT.n4 OUT.n26 0.042
R120 OUT.n3 OUT.n17 0.042
R121 OUT.n2 OUT.n20 0.042
R122 OUT.n1 OUT.n11 0.042
R123 OUT.n0 OUT.n7 0.042
R124 OUT.n6 OUT.n5 0.039
R125 OUT.n10 OUT.n9 0.039
R126 OUT.n16 OUT.n15 0.039
R127 OUT.n25 OUT.n24 0.039
R128 VDD.n13 VDD.n12 101.754
R129 VDD.n22 VDD.n0 99.531
R130 VDD.n6 VDD.n4 99.225
R131 VDD.n24 VDD.n23 96.689
R132 VDD.n6 VDD.n5 96.506
R133 VDD.n22 VDD.n14 96.445
R134 VDD.n26 VDD.n25 96.383
R135 VDD.n3 VDD.n1 96.199
R136 VDD.n9 VDD.n8 96.077
R137 VDD.n28 VDD.n27 96.016
R138 VDD.n3 VDD.n2 19.259
R139 VDD.n12 VDD.t6 8
R140 VDD.n8 VDD.t7 7.998
R141 VDD.n1 VDD.t4 7.998
R142 VDD.n14 VDD.t19 7.998
R143 VDD.n23 VDD.t18 7.998
R144 VDD.n27 VDD.t15 7.998
R145 VDD.n25 VDD.t17 7.998
R146 VDD.n4 VDD.t0 7.998
R147 VDD.n5 VDD.t9 7.998
R148 VDD.n21 VDD.t16 7.917
R149 VDD.n8 VDD.t8 6.181
R150 VDD.n1 VDD.t3 6.181
R151 VDD.n14 VDD.t13 6.181
R152 VDD.n23 VDD.t11 6.181
R153 VDD.n27 VDD.t12 6.181
R154 VDD.n25 VDD.t10 6.181
R155 VDD.n4 VDD.t2 6.181
R156 VDD.n5 VDD.t5 6.181
R157 VDD.n12 VDD.t1 6.173
R158 VDD.n15 VDD.t14 5.809
R159 VDD.n10 VDD.n9 0.362
R160 VDD VDD.n28 0.271
R161 VDD VDD.n13 0.262
R162 VDD.n24 VDD.n22 0.189
R163 VDD.n10 VDD.n7 0.189
R164 VDD.n26 VDD.n24 0.188
R165 VDD.n7 VDD.n6 0.187
R166 VDD.n7 VDD.n3 0.185
R167 VDD.n28 VDD.n26 0.178
R168 VDD.n13 VDD.n11 0.14
R169 VDD.n0 VDD.n20 0.083
R170 VDD.n0 VDD.n21 0.082
R171 VDD.n16 VDD.n15 0.082
R172 VDD.n18 VDD.n17 0.082
R173 VDD.n20 VDD.n19 0.06
R174 VDD.n17 VDD.n16 0.041
R175 VDD.n11 VDD.n10 0.038
R176 VDD.n19 VDD.n18 0.023
R177 GND.n1 GND.t3 78.958
R178 GND.n3 GND.n2 56.838
R179 GND.n1 GND.n0 56.822
R180 GND.n2 GND.t1 25.253
R181 GND.n2 GND.t2 24.558
R182 GND.n0 GND.t4 24.418
R183 GND.n0 GND.t0 24.137
R184 GND GND.n3 0.639
R185 GND.n3 GND.n1 0.434
C0 A w_n15748_5772# 0.41fF
C1 IN GND 1.13fF
C2 VDD w_n15748_5772# 0.25fF
C3 OUT w_n3748_5772# 0.41fF
C4 OUT IN 0.79fF
C5 OUT A 1.24fF
C6 w_n3748_5772# VDD 0.25fF
C7 GND VSUBS 10.78fF $ **FLOATING
C8 IN VSUBS 11.75fF
C9 OUT VSUBS 16.07fF $ **FLOATING
C10 VDD VSUBS 43.96fF $ **FLOATING
C11 A VSUBS 62.77fF $ **FLOATING
C12 w_n3748_5772# VSUBS 315.49fF
C13 w_n15748_5772# VSUBS 315.49fF
C14 GND.t4 VSUBS 0.28fF
C15 GND.t0 VSUBS 0.27fF
C16 GND.n0 VSUBS 0.78fF $ **FLOATING
C17 GND.t3 VSUBS 0.91fF
C18 GND.n1 VSUBS 2.28fF $ **FLOATING
C19 GND.t2 VSUBS 0.28fF
C20 GND.t1 VSUBS 0.29fF
C21 GND.n2 VSUBS 0.76fF $ **FLOATING
C22 GND.n3 VSUBS 1.33fF $ **FLOATING
C23 VDD.n0 VSUBS 0.15fF $ **FLOATING
C24 VDD.t4 VSUBS 0.68fF
C25 VDD.t3 VSUBS 0.54fF
C26 VDD.n1 VSUBS 1.93fF $ **FLOATING
C27 VDD.n2 VSUBS 0.17fF $ **FLOATING
C28 VDD.n3 VSUBS 0.10fF $ **FLOATING
C29 VDD.t0 VSUBS 0.68fF
C30 VDD.t2 VSUBS 0.54fF
C31 VDD.n4 VSUBS 1.93fF $ **FLOATING
C32 VDD.t9 VSUBS 0.68fF
C33 VDD.t5 VSUBS 0.54fF
C34 VDD.n5 VSUBS 1.93fF $ **FLOATING
C35 VDD.n6 VSUBS 1.95fF $ **FLOATING
C36 VDD.n7 VSUBS 0.90fF $ **FLOATING
C37 VDD.t7 VSUBS 0.68fF
C38 VDD.t8 VSUBS 0.54fF
C39 VDD.n8 VSUBS 1.93fF $ **FLOATING
C40 VDD.n9 VSUBS 0.10fF $ **FLOATING
C41 VDD.n10 VSUBS 0.76fF $ **FLOATING
C42 VDD.n11 VSUBS 0.19fF $ **FLOATING
C43 VDD.t6 VSUBS 0.68fF
C44 VDD.t1 VSUBS 0.26fF
C45 VDD.n12 VSUBS 2.21fF $ **FLOATING
C46 VDD.n13 VSUBS 1.01fF $ **FLOATING
C47 VDD.t19 VSUBS 0.68fF
C48 VDD.t13 VSUBS 0.54fF
C49 VDD.n14 VSUBS 1.93fF $ **FLOATING
C50 VDD.t14 VSUBS 0.19fF
C51 VDD.n15 VSUBS 0.86fF $ **FLOATING
C52 VDD.n16 VSUBS 0.11fF $ **FLOATING
C53 VDD.n17 VSUBS 0.08fF $ **FLOATING
C54 VDD.n18 VSUBS 0.18fF $ **FLOATING
C55 VDD.n20 VSUBS 0.18fF $ **FLOATING
C56 VDD.t16 VSUBS 0.67fF
C57 VDD.n21 VSUBS 0.74fF $ **FLOATING
C58 VDD.n22 VSUBS 1.86fF $ **FLOATING
C59 VDD.t18 VSUBS 0.68fF
C60 VDD.t11 VSUBS 0.54fF
C61 VDD.n23 VSUBS 1.93fF $ **FLOATING
C62 VDD.n24 VSUBS 1.07fF $ **FLOATING
C63 VDD.t17 VSUBS 0.68fF
C64 VDD.t10 VSUBS 0.54fF
C65 VDD.n25 VSUBS 1.93fF $ **FLOATING
C66 VDD.n26 VSUBS 1.05fF $ **FLOATING
C67 VDD.t15 VSUBS 0.68fF
C68 VDD.t12 VSUBS 0.54fF
C69 VDD.n27 VSUBS 1.93fF $ **FLOATING
C70 VDD.n28 VSUBS 1.13fF $ **FLOATING
C71 OUT.n0 VSUBS 0.07fF $ **FLOATING
C72 OUT.n1 VSUBS 0.07fF $ **FLOATING
C73 OUT.n2 VSUBS 0.25fF $ **FLOATING
C74 OUT.n3 VSUBS 0.07fF $ **FLOATING
C75 OUT.n4 VSUBS 0.07fF $ **FLOATING
C76 OUT.t12 VSUBS 0.35fF
C77 OUT.n5 VSUBS 0.40fF $ **FLOATING
C78 OUT.n7 VSUBS 0.08fF $ **FLOATING
C79 OUT.n8 VSUBS 0.83fF $ **FLOATING
C80 OUT.t7 VSUBS 0.35fF
C81 OUT.n9 VSUBS 0.40fF $ **FLOATING
C82 OUT.n11 VSUBS 0.08fF $ **FLOATING
C83 OUT.n12 VSUBS 0.83fF $ **FLOATING
C84 OUT.t14 VSUBS 1.42fF
C85 OUT.n13 VSUBS 0.67fF $ **FLOATING
C86 OUT.n14 VSUBS 0.11fF $ **FLOATING
C87 OUT.t8 VSUBS 0.35fF
C88 OUT.n15 VSUBS 0.40fF $ **FLOATING
C89 OUT.n17 VSUBS 0.08fF $ **FLOATING
C90 OUT.n18 VSUBS 0.83fF $ **FLOATING
C91 OUT.n20 VSUBS 1.36fF $ **FLOATING
C92 OUT.t13 VSUBS 0.48fF
C93 OUT.n21 VSUBS 0.53fF $ **FLOATING
C94 OUT.n22 VSUBS 0.20fF $ **FLOATING
C95 OUT.n23 VSUBS 0.18fF $ **FLOATING
C96 OUT.t5 VSUBS 0.35fF
C97 OUT.n24 VSUBS 0.40fF $ **FLOATING
C98 OUT.n26 VSUBS 0.08fF $ **FLOATING
C99 OUT.n27 VSUBS 0.83fF $ **FLOATING
C100 OUT.n28 VSUBS 0.11fF $ **FLOATING
C101 OUT.n29 VSUBS 0.09fF $ **FLOATING
C102 OUT.t2 VSUBS 0.35fF
C103 OUT.t1 VSUBS 0.07fF
C104 OUT.t0 VSUBS 0.06fF
C105 OUT.n30 VSUBS 0.23fF $ **FLOATING
C106 OUT.t3 VSUBS 0.07fF
C107 OUT.t4 VSUBS 0.08fF
C108 OUT.n31 VSUBS 0.21fF $ **FLOATING
C109 OUT.n32 VSUBS 0.26fF $ **FLOATING
C110 OUT.t6 VSUBS 0.50fF
C111 OUT.t10 VSUBS 0.50fF
C112 OUT.t11 VSUBS 0.50fF
C113 OUT.t9 VSUBS 0.50fF
C114 A.n0 VSUBS 0.49fF $ **FLOATING
C115 A.n1 VSUBS 0.17fF $ **FLOATING
C116 A.n2 VSUBS 0.17fF $ **FLOATING
C117 A.n3 VSUBS 0.17fF $ **FLOATING
C118 A.n4 VSUBS 0.17fF $ **FLOATING
C119 A.t8 VSUBS 0.87fF
C120 A.t10 VSUBS 0.87fF
C121 A.t6 VSUBS 0.87fF
C122 A.t4 VSUBS 0.87fF
C123 A.t12 VSUBS 0.87fF
C124 A.t16 VSUBS 0.87fF
C125 A.t14 VSUBS 0.87fF
C126 A.t0 VSUBS 0.87fF
C127 A.t18 VSUBS 0.87fF
C128 A.t2 VSUBS 0.93fF
C129 A.n5 VSUBS 0.81fF $ **FLOATING
C130 A.n6 VSUBS 0.46fF $ **FLOATING
C131 A.n7 VSUBS 0.46fF $ **FLOATING
C132 A.n8 VSUBS 0.46fF $ **FLOATING
C133 A.n9 VSUBS 0.46fF $ **FLOATING
C134 A.n10 VSUBS 0.46fF $ **FLOATING
C135 A.n11 VSUBS 0.46fF $ **FLOATING
C136 A.n12 VSUBS 0.46fF $ **FLOATING
C137 A.n13 VSUBS 0.53fF $ **FLOATING
C138 A.t23 VSUBS 0.87fF
C139 A.t28 VSUBS 0.87fF
C140 A.t22 VSUBS 0.87fF
C141 A.t21 VSUBS 0.87fF
C142 A.t25 VSUBS 0.87fF
C143 A.t26 VSUBS 0.87fF
C144 A.t20 VSUBS 0.87fF
C145 A.t24 VSUBS 0.87fF
C146 A.t29 VSUBS 0.87fF
C147 A.t27 VSUBS 0.93fF
C148 A.n14 VSUBS 0.81fF $ **FLOATING
C149 A.n15 VSUBS 0.46fF $ **FLOATING
C150 A.n16 VSUBS 0.46fF $ **FLOATING
C151 A.n17 VSUBS 0.46fF $ **FLOATING
C152 A.n18 VSUBS 0.46fF $ **FLOATING
C153 A.n19 VSUBS 0.46fF $ **FLOATING
C154 A.n20 VSUBS 0.46fF $ **FLOATING
C155 A.n21 VSUBS 0.46fF $ **FLOATING
C156 A.n22 VSUBS 0.50fF $ **FLOATING
C157 A.n23 VSUBS 0.70fF $ **FLOATING
C158 A.n24 VSUBS 0.01fF $ **FLOATING
C159 A.n25 VSUBS 3.32fF $ **FLOATING
C160 A.t9 VSUBS 1.17fF
C161 A.n26 VSUBS 1.29fF $ **FLOATING
C162 A.n27 VSUBS 0.48fF $ **FLOATING
C163 A.t11 VSUBS 0.86fF
C164 A.n28 VSUBS 0.97fF $ **FLOATING
C165 A.n30 VSUBS 0.18fF $ **FLOATING
C166 A.n31 VSUBS 2.04fF $ **FLOATING
C167 A.t5 VSUBS 0.86fF
C168 A.n32 VSUBS 0.97fF $ **FLOATING
C169 A.n34 VSUBS 0.18fF $ **FLOATING
C170 A.n35 VSUBS 2.04fF $ **FLOATING
C171 A.t17 VSUBS 0.86fF
C172 A.n36 VSUBS 0.97fF $ **FLOATING
C173 A.n38 VSUBS 0.18fF $ **FLOATING
C174 A.n39 VSUBS 2.04fF $ **FLOATING
C175 A.t3 VSUBS 3.47fF
C176 A.t1 VSUBS 0.86fF
C177 A.n40 VSUBS 0.97fF $ **FLOATING
C178 A.n42 VSUBS 0.18fF $ **FLOATING
C179 A.n43 VSUBS 2.04fF $ **FLOATING
C180 A.n44 VSUBS 1.63fF $ **FLOATING
C181 A.n45 VSUBS 0.33fF $ **FLOATING
C182 A.n46 VSUBS 0.34fF $ **FLOATING
C183 A.n47 VSUBS 0.33fF $ **FLOATING
C184 A.n48 VSUBS 0.32fF $ **FLOATING
C185 A.n49 VSUBS 0.34fF $ **FLOATING
C186 A.t7 VSUBS 1.22fF
C187 A.t13 VSUBS 1.22fF
C188 A.t15 VSUBS 1.22fF
C189 A.t19 VSUBS 1.22fF
.ends
