magic
tech sky130A
timestamp 1621261496
<< nwell >>
rect -7874 2886 -2726 7970
rect -1874 2886 3274 7970
rect -7764 2863 -2726 2886
rect -1764 2863 3274 2886
rect -7237 2862 -6570 2863
rect -6347 2862 -6125 2863
rect -5902 2862 -5680 2863
rect -5457 2862 -5235 2863
rect -5012 2862 -4790 2863
rect -4567 2862 -4345 2863
rect -4122 2862 -3900 2863
rect -3677 2862 -3455 2863
rect -3232 2862 -3010 2863
rect -1237 2862 -570 2863
rect -347 2862 -125 2863
rect 98 2862 320 2863
rect 543 2862 765 2863
rect 988 2862 1210 2863
rect 1433 2862 1655 2863
rect 1878 2862 2100 2863
rect 2323 2862 2545 2863
rect 2768 2862 2990 2863
<< nmos >>
rect 0 -13 100 847
rect 457 -13 557 847
rect 905 -13 1005 847
rect 1353 -13 1453 847
rect 1746 -13 1846 847
<< pmos >>
rect -7460 3047 -7360 7837
rect -7015 3046 -6915 7837
rect -6570 3046 -6470 7837
rect -6125 3046 -6025 7837
rect -5680 3046 -5580 7837
rect -5235 3046 -5135 7837
rect -4790 3046 -4690 7837
rect -4345 3046 -4245 7837
rect -3900 3046 -3800 7837
rect -3455 3046 -3355 7837
rect -1460 3047 -1360 7837
rect -1015 3046 -915 7837
rect -570 3046 -470 7837
rect -125 3046 -25 7837
rect 320 3046 420 7837
rect 765 3046 865 7837
rect 1210 3046 1310 7837
rect 1655 3046 1755 7837
rect 2100 3046 2200 7837
rect 2545 3046 2645 7837
<< ndiff >>
rect -329 606 0 847
rect -329 506 -232 606
rect -132 506 0 606
rect -329 373 0 506
rect -329 273 -234 373
rect -134 273 0 373
rect -329 -13 0 273
rect 100 606 457 847
rect 100 506 228 606
rect 328 506 457 606
rect 100 373 457 506
rect 100 273 226 373
rect 326 273 457 373
rect 100 -13 457 273
rect 557 608 905 847
rect 557 508 668 608
rect 768 508 905 608
rect 557 375 905 508
rect 557 275 666 375
rect 766 275 905 375
rect 557 -13 905 275
rect 1005 608 1353 847
rect 1005 508 1132 608
rect 1232 508 1353 608
rect 1005 375 1353 508
rect 1005 275 1130 375
rect 1230 275 1353 375
rect 1005 -13 1353 275
rect 1453 610 1746 847
rect 1453 510 1558 610
rect 1658 510 1746 610
rect 1453 377 1746 510
rect 1453 277 1556 377
rect 1656 277 1746 377
rect 1453 -13 1746 277
rect 1846 610 2148 847
rect 1846 510 1953 610
rect 2053 510 2148 610
rect 1846 377 2148 510
rect 1846 277 1951 377
rect 2051 277 2148 377
rect 1846 -13 2148 277
<< pdiff >>
rect -7730 7778 -7460 7837
rect -7730 7707 -7628 7778
rect -7557 7707 -7460 7778
rect -7730 7459 -7460 7707
rect -7730 7388 -7624 7459
rect -7553 7388 -7460 7459
rect -7730 7133 -7460 7388
rect -7730 7062 -7621 7133
rect -7550 7062 -7460 7133
rect -7730 6882 -7460 7062
rect -7730 6811 -7624 6882
rect -7553 6811 -7460 6882
rect -7730 6604 -7460 6811
rect -7730 6533 -7624 6604
rect -7553 6533 -7460 6604
rect -7730 6353 -7460 6533
rect -7730 6282 -7624 6353
rect -7553 6282 -7460 6353
rect -7730 6031 -7460 6282
rect -7730 5960 -7628 6031
rect -7557 5960 -7460 6031
rect -7730 5690 -7460 5960
rect -7730 5619 -7621 5690
rect -7550 5619 -7460 5690
rect -7730 5307 -7460 5619
rect -7730 5236 -7626 5307
rect -7555 5236 -7460 5307
rect -7730 4945 -7460 5236
rect -7730 4874 -7626 4945
rect -7555 4874 -7460 4945
rect -7730 4602 -7460 4874
rect -7730 4531 -7619 4602
rect -7548 4531 -7460 4602
rect -7730 4184 -7460 4531
rect -7730 4113 -7630 4184
rect -7559 4113 -7460 4184
rect -7730 3769 -7460 4113
rect -7730 3698 -7626 3769
rect -7555 3698 -7460 3769
rect -7730 3399 -7460 3698
rect -7730 3328 -7622 3399
rect -7551 3328 -7460 3399
rect -7730 3047 -7460 3328
rect -7360 7777 -7015 7837
rect -7360 7706 -7201 7777
rect -7130 7706 -7015 7777
rect -7360 7458 -7015 7706
rect -7360 7387 -7197 7458
rect -7126 7387 -7015 7458
rect -7360 7132 -7015 7387
rect -7360 7061 -7194 7132
rect -7123 7061 -7015 7132
rect -7360 6881 -7015 7061
rect -7360 6810 -7197 6881
rect -7126 6810 -7015 6881
rect -7360 6603 -7015 6810
rect -7360 6532 -7197 6603
rect -7126 6532 -7015 6603
rect -7360 6352 -7015 6532
rect -7360 6281 -7197 6352
rect -7126 6281 -7015 6352
rect -7360 6030 -7015 6281
rect -7360 5959 -7201 6030
rect -7130 5959 -7015 6030
rect -7360 5689 -7015 5959
rect -7360 5618 -7194 5689
rect -7123 5618 -7015 5689
rect -7360 5306 -7015 5618
rect -7360 5235 -7199 5306
rect -7128 5235 -7015 5306
rect -7360 4944 -7015 5235
rect -7360 4873 -7199 4944
rect -7128 4873 -7015 4944
rect -7360 4601 -7015 4873
rect -7360 4530 -7192 4601
rect -7121 4530 -7015 4601
rect -7360 4183 -7015 4530
rect -7360 4112 -7203 4183
rect -7132 4112 -7015 4183
rect -7360 3768 -7015 4112
rect -7360 3697 -7199 3768
rect -7128 3697 -7015 3768
rect -7360 3398 -7015 3697
rect -7360 3327 -7195 3398
rect -7124 3327 -7015 3398
rect -7360 3047 -7015 3327
rect -7237 3046 -7015 3047
rect -6915 7777 -6570 7837
rect -6915 7706 -6756 7777
rect -6685 7706 -6570 7777
rect -6915 7458 -6570 7706
rect -6915 7387 -6752 7458
rect -6681 7387 -6570 7458
rect -6915 7132 -6570 7387
rect -6915 7061 -6749 7132
rect -6678 7061 -6570 7132
rect -6915 6881 -6570 7061
rect -6915 6810 -6752 6881
rect -6681 6810 -6570 6881
rect -6915 6603 -6570 6810
rect -6915 6532 -6752 6603
rect -6681 6532 -6570 6603
rect -6915 6352 -6570 6532
rect -6915 6281 -6752 6352
rect -6681 6281 -6570 6352
rect -6915 6030 -6570 6281
rect -6915 5959 -6756 6030
rect -6685 5959 -6570 6030
rect -6915 5689 -6570 5959
rect -6915 5618 -6749 5689
rect -6678 5618 -6570 5689
rect -6915 5306 -6570 5618
rect -6915 5235 -6754 5306
rect -6683 5235 -6570 5306
rect -6915 4944 -6570 5235
rect -6915 4873 -6754 4944
rect -6683 4873 -6570 4944
rect -6915 4601 -6570 4873
rect -6915 4530 -6747 4601
rect -6676 4530 -6570 4601
rect -6915 4183 -6570 4530
rect -6915 4112 -6758 4183
rect -6687 4112 -6570 4183
rect -6915 3768 -6570 4112
rect -6915 3697 -6754 3768
rect -6683 3697 -6570 3768
rect -6915 3398 -6570 3697
rect -6915 3327 -6750 3398
rect -6679 3327 -6570 3398
rect -6915 3046 -6570 3327
rect -6470 7777 -6125 7837
rect -6470 7706 -6311 7777
rect -6240 7706 -6125 7777
rect -6470 7458 -6125 7706
rect -6470 7387 -6307 7458
rect -6236 7387 -6125 7458
rect -6470 7132 -6125 7387
rect -6470 7061 -6304 7132
rect -6233 7061 -6125 7132
rect -6470 6881 -6125 7061
rect -6470 6810 -6307 6881
rect -6236 6810 -6125 6881
rect -6470 6603 -6125 6810
rect -6470 6532 -6307 6603
rect -6236 6532 -6125 6603
rect -6470 6352 -6125 6532
rect -6470 6281 -6307 6352
rect -6236 6281 -6125 6352
rect -6470 6030 -6125 6281
rect -6470 5959 -6311 6030
rect -6240 5959 -6125 6030
rect -6470 5689 -6125 5959
rect -6470 5618 -6304 5689
rect -6233 5618 -6125 5689
rect -6470 5306 -6125 5618
rect -6470 5235 -6309 5306
rect -6238 5235 -6125 5306
rect -6470 4944 -6125 5235
rect -6470 4873 -6309 4944
rect -6238 4873 -6125 4944
rect -6470 4601 -6125 4873
rect -6470 4530 -6302 4601
rect -6231 4530 -6125 4601
rect -6470 4183 -6125 4530
rect -6470 4112 -6313 4183
rect -6242 4112 -6125 4183
rect -6470 3768 -6125 4112
rect -6470 3697 -6309 3768
rect -6238 3697 -6125 3768
rect -6470 3398 -6125 3697
rect -6470 3327 -6305 3398
rect -6234 3327 -6125 3398
rect -6470 3046 -6125 3327
rect -6025 7777 -5680 7837
rect -6025 7706 -5866 7777
rect -5795 7706 -5680 7777
rect -6025 7458 -5680 7706
rect -6025 7387 -5862 7458
rect -5791 7387 -5680 7458
rect -6025 7132 -5680 7387
rect -6025 7061 -5859 7132
rect -5788 7061 -5680 7132
rect -6025 6881 -5680 7061
rect -6025 6810 -5862 6881
rect -5791 6810 -5680 6881
rect -6025 6603 -5680 6810
rect -6025 6532 -5862 6603
rect -5791 6532 -5680 6603
rect -6025 6352 -5680 6532
rect -6025 6281 -5862 6352
rect -5791 6281 -5680 6352
rect -6025 6030 -5680 6281
rect -6025 5959 -5866 6030
rect -5795 5959 -5680 6030
rect -6025 5689 -5680 5959
rect -6025 5618 -5859 5689
rect -5788 5618 -5680 5689
rect -6025 5306 -5680 5618
rect -6025 5235 -5864 5306
rect -5793 5235 -5680 5306
rect -6025 4944 -5680 5235
rect -6025 4873 -5864 4944
rect -5793 4873 -5680 4944
rect -6025 4601 -5680 4873
rect -6025 4530 -5857 4601
rect -5786 4530 -5680 4601
rect -6025 4183 -5680 4530
rect -6025 4112 -5868 4183
rect -5797 4112 -5680 4183
rect -6025 3768 -5680 4112
rect -6025 3697 -5864 3768
rect -5793 3697 -5680 3768
rect -6025 3398 -5680 3697
rect -6025 3327 -5860 3398
rect -5789 3327 -5680 3398
rect -6025 3046 -5680 3327
rect -5580 7777 -5235 7837
rect -5580 7706 -5421 7777
rect -5350 7706 -5235 7777
rect -5580 7458 -5235 7706
rect -5580 7387 -5417 7458
rect -5346 7387 -5235 7458
rect -5580 7132 -5235 7387
rect -5580 7061 -5414 7132
rect -5343 7061 -5235 7132
rect -5580 6881 -5235 7061
rect -5580 6810 -5417 6881
rect -5346 6810 -5235 6881
rect -5580 6603 -5235 6810
rect -5580 6532 -5417 6603
rect -5346 6532 -5235 6603
rect -5580 6352 -5235 6532
rect -5580 6281 -5417 6352
rect -5346 6281 -5235 6352
rect -5580 6030 -5235 6281
rect -5580 5959 -5421 6030
rect -5350 5959 -5235 6030
rect -5580 5689 -5235 5959
rect -5580 5618 -5414 5689
rect -5343 5618 -5235 5689
rect -5580 5306 -5235 5618
rect -5580 5235 -5419 5306
rect -5348 5235 -5235 5306
rect -5580 4944 -5235 5235
rect -5580 4873 -5419 4944
rect -5348 4873 -5235 4944
rect -5580 4601 -5235 4873
rect -5580 4530 -5412 4601
rect -5341 4530 -5235 4601
rect -5580 4183 -5235 4530
rect -5580 4112 -5423 4183
rect -5352 4112 -5235 4183
rect -5580 3768 -5235 4112
rect -5580 3697 -5419 3768
rect -5348 3697 -5235 3768
rect -5580 3398 -5235 3697
rect -5580 3327 -5415 3398
rect -5344 3327 -5235 3398
rect -5580 3046 -5235 3327
rect -5135 7777 -4790 7837
rect -5135 7706 -4976 7777
rect -4905 7706 -4790 7777
rect -5135 7458 -4790 7706
rect -5135 7387 -4972 7458
rect -4901 7387 -4790 7458
rect -5135 7132 -4790 7387
rect -5135 7061 -4969 7132
rect -4898 7061 -4790 7132
rect -5135 6881 -4790 7061
rect -5135 6810 -4972 6881
rect -4901 6810 -4790 6881
rect -5135 6603 -4790 6810
rect -5135 6532 -4972 6603
rect -4901 6532 -4790 6603
rect -5135 6352 -4790 6532
rect -5135 6281 -4972 6352
rect -4901 6281 -4790 6352
rect -5135 6030 -4790 6281
rect -5135 5959 -4976 6030
rect -4905 5959 -4790 6030
rect -5135 5689 -4790 5959
rect -5135 5618 -4969 5689
rect -4898 5618 -4790 5689
rect -5135 5306 -4790 5618
rect -5135 5235 -4974 5306
rect -4903 5235 -4790 5306
rect -5135 4944 -4790 5235
rect -5135 4873 -4974 4944
rect -4903 4873 -4790 4944
rect -5135 4601 -4790 4873
rect -5135 4530 -4967 4601
rect -4896 4530 -4790 4601
rect -5135 4183 -4790 4530
rect -5135 4112 -4978 4183
rect -4907 4112 -4790 4183
rect -5135 3768 -4790 4112
rect -5135 3697 -4974 3768
rect -4903 3697 -4790 3768
rect -5135 3398 -4790 3697
rect -5135 3327 -4970 3398
rect -4899 3327 -4790 3398
rect -5135 3046 -4790 3327
rect -4690 7777 -4345 7837
rect -4690 7706 -4531 7777
rect -4460 7706 -4345 7777
rect -4690 7458 -4345 7706
rect -4690 7387 -4527 7458
rect -4456 7387 -4345 7458
rect -4690 7132 -4345 7387
rect -4690 7061 -4524 7132
rect -4453 7061 -4345 7132
rect -4690 6881 -4345 7061
rect -4690 6810 -4527 6881
rect -4456 6810 -4345 6881
rect -4690 6603 -4345 6810
rect -4690 6532 -4527 6603
rect -4456 6532 -4345 6603
rect -4690 6352 -4345 6532
rect -4690 6281 -4527 6352
rect -4456 6281 -4345 6352
rect -4690 6030 -4345 6281
rect -4690 5959 -4531 6030
rect -4460 5959 -4345 6030
rect -4690 5689 -4345 5959
rect -4690 5618 -4524 5689
rect -4453 5618 -4345 5689
rect -4690 5306 -4345 5618
rect -4690 5235 -4529 5306
rect -4458 5235 -4345 5306
rect -4690 4944 -4345 5235
rect -4690 4873 -4529 4944
rect -4458 4873 -4345 4944
rect -4690 4601 -4345 4873
rect -4690 4530 -4522 4601
rect -4451 4530 -4345 4601
rect -4690 4183 -4345 4530
rect -4690 4112 -4533 4183
rect -4462 4112 -4345 4183
rect -4690 3768 -4345 4112
rect -4690 3697 -4529 3768
rect -4458 3697 -4345 3768
rect -4690 3398 -4345 3697
rect -4690 3327 -4525 3398
rect -4454 3327 -4345 3398
rect -4690 3046 -4345 3327
rect -4245 7777 -3900 7837
rect -4245 7706 -4086 7777
rect -4015 7706 -3900 7777
rect -4245 7458 -3900 7706
rect -4245 7387 -4082 7458
rect -4011 7387 -3900 7458
rect -4245 7132 -3900 7387
rect -4245 7061 -4079 7132
rect -4008 7061 -3900 7132
rect -4245 6881 -3900 7061
rect -4245 6810 -4082 6881
rect -4011 6810 -3900 6881
rect -4245 6603 -3900 6810
rect -4245 6532 -4082 6603
rect -4011 6532 -3900 6603
rect -4245 6352 -3900 6532
rect -4245 6281 -4082 6352
rect -4011 6281 -3900 6352
rect -4245 6030 -3900 6281
rect -4245 5959 -4086 6030
rect -4015 5959 -3900 6030
rect -4245 5689 -3900 5959
rect -4245 5618 -4079 5689
rect -4008 5618 -3900 5689
rect -4245 5306 -3900 5618
rect -4245 5235 -4084 5306
rect -4013 5235 -3900 5306
rect -4245 4944 -3900 5235
rect -4245 4873 -4084 4944
rect -4013 4873 -3900 4944
rect -4245 4601 -3900 4873
rect -4245 4530 -4077 4601
rect -4006 4530 -3900 4601
rect -4245 4183 -3900 4530
rect -4245 4112 -4088 4183
rect -4017 4112 -3900 4183
rect -4245 3768 -3900 4112
rect -4245 3697 -4084 3768
rect -4013 3697 -3900 3768
rect -4245 3398 -3900 3697
rect -4245 3327 -4080 3398
rect -4009 3327 -3900 3398
rect -4245 3046 -3900 3327
rect -3800 7777 -3455 7837
rect -3800 7706 -3641 7777
rect -3570 7706 -3455 7777
rect -3800 7458 -3455 7706
rect -3800 7387 -3637 7458
rect -3566 7387 -3455 7458
rect -3800 7132 -3455 7387
rect -3800 7061 -3634 7132
rect -3563 7061 -3455 7132
rect -3800 6881 -3455 7061
rect -3800 6810 -3637 6881
rect -3566 6810 -3455 6881
rect -3800 6603 -3455 6810
rect -3800 6532 -3637 6603
rect -3566 6532 -3455 6603
rect -3800 6352 -3455 6532
rect -3800 6281 -3637 6352
rect -3566 6281 -3455 6352
rect -3800 6030 -3455 6281
rect -3800 5959 -3641 6030
rect -3570 5959 -3455 6030
rect -3800 5689 -3455 5959
rect -3800 5618 -3634 5689
rect -3563 5618 -3455 5689
rect -3800 5306 -3455 5618
rect -3800 5235 -3639 5306
rect -3568 5235 -3455 5306
rect -3800 4944 -3455 5235
rect -3800 4873 -3639 4944
rect -3568 4873 -3455 4944
rect -3800 4601 -3455 4873
rect -3800 4530 -3632 4601
rect -3561 4530 -3455 4601
rect -3800 4183 -3455 4530
rect -3800 4112 -3643 4183
rect -3572 4112 -3455 4183
rect -3800 3768 -3455 4112
rect -3800 3697 -3639 3768
rect -3568 3697 -3455 3768
rect -3800 3398 -3455 3697
rect -3800 3327 -3635 3398
rect -3564 3327 -3455 3398
rect -3800 3046 -3455 3327
rect -3355 7777 -2902 7837
rect -3355 7706 -3196 7777
rect -3125 7706 -2902 7777
rect -3355 7458 -2902 7706
rect -3355 7387 -3192 7458
rect -3121 7387 -2902 7458
rect -3355 7132 -2902 7387
rect -3355 7061 -3189 7132
rect -3118 7061 -2902 7132
rect -3355 6881 -2902 7061
rect -3355 6810 -3192 6881
rect -3121 6810 -2902 6881
rect -3355 6603 -2902 6810
rect -3355 6532 -3192 6603
rect -3121 6532 -2902 6603
rect -3355 6352 -2902 6532
rect -3355 6281 -3192 6352
rect -3121 6281 -2902 6352
rect -3355 6030 -2902 6281
rect -3355 5959 -3196 6030
rect -3125 5959 -2902 6030
rect -3355 5689 -2902 5959
rect -3355 5618 -3189 5689
rect -3118 5618 -2902 5689
rect -3355 5306 -2902 5618
rect -3355 5235 -3194 5306
rect -3123 5235 -2902 5306
rect -3355 4944 -2902 5235
rect -3355 4873 -3194 4944
rect -3123 4873 -2902 4944
rect -3355 4601 -2902 4873
rect -3355 4530 -3187 4601
rect -3116 4530 -2902 4601
rect -3355 4183 -2902 4530
rect -3355 4112 -3198 4183
rect -3127 4112 -2902 4183
rect -3355 3768 -2902 4112
rect -3355 3697 -3194 3768
rect -3123 3697 -2902 3768
rect -3355 3398 -2902 3697
rect -3355 3327 -3190 3398
rect -3119 3327 -2902 3398
rect -3355 3062 -2902 3327
rect -1730 7778 -1460 7837
rect -1730 7707 -1628 7778
rect -1557 7707 -1460 7778
rect -1730 7459 -1460 7707
rect -1730 7388 -1624 7459
rect -1553 7388 -1460 7459
rect -1730 7133 -1460 7388
rect -1730 7062 -1621 7133
rect -1550 7062 -1460 7133
rect -1730 6882 -1460 7062
rect -1730 6811 -1624 6882
rect -1553 6811 -1460 6882
rect -1730 6604 -1460 6811
rect -1730 6533 -1624 6604
rect -1553 6533 -1460 6604
rect -1730 6353 -1460 6533
rect -1730 6282 -1624 6353
rect -1553 6282 -1460 6353
rect -1730 6031 -1460 6282
rect -1730 5960 -1628 6031
rect -1557 5960 -1460 6031
rect -1730 5690 -1460 5960
rect -1730 5619 -1621 5690
rect -1550 5619 -1460 5690
rect -1730 5307 -1460 5619
rect -1730 5236 -1626 5307
rect -1555 5236 -1460 5307
rect -1730 4945 -1460 5236
rect -1730 4874 -1626 4945
rect -1555 4874 -1460 4945
rect -1730 4602 -1460 4874
rect -1730 4531 -1619 4602
rect -1548 4531 -1460 4602
rect -1730 4184 -1460 4531
rect -1730 4113 -1630 4184
rect -1559 4113 -1460 4184
rect -1730 3769 -1460 4113
rect -1730 3698 -1626 3769
rect -1555 3698 -1460 3769
rect -1730 3399 -1460 3698
rect -1730 3328 -1622 3399
rect -1551 3328 -1460 3399
rect -3355 3046 -2901 3062
rect -1730 3047 -1460 3328
rect -1360 7777 -1015 7837
rect -1360 7706 -1201 7777
rect -1130 7706 -1015 7777
rect -1360 7458 -1015 7706
rect -1360 7387 -1197 7458
rect -1126 7387 -1015 7458
rect -1360 7132 -1015 7387
rect -1360 7061 -1194 7132
rect -1123 7061 -1015 7132
rect -1360 6881 -1015 7061
rect -1360 6810 -1197 6881
rect -1126 6810 -1015 6881
rect -1360 6603 -1015 6810
rect -1360 6532 -1197 6603
rect -1126 6532 -1015 6603
rect -1360 6352 -1015 6532
rect -1360 6281 -1197 6352
rect -1126 6281 -1015 6352
rect -1360 6030 -1015 6281
rect -1360 5959 -1201 6030
rect -1130 5959 -1015 6030
rect -1360 5689 -1015 5959
rect -1360 5618 -1194 5689
rect -1123 5618 -1015 5689
rect -1360 5306 -1015 5618
rect -1360 5235 -1199 5306
rect -1128 5235 -1015 5306
rect -1360 4944 -1015 5235
rect -1360 4873 -1199 4944
rect -1128 4873 -1015 4944
rect -1360 4601 -1015 4873
rect -1360 4530 -1192 4601
rect -1121 4530 -1015 4601
rect -1360 4183 -1015 4530
rect -1360 4112 -1203 4183
rect -1132 4112 -1015 4183
rect -1360 3768 -1015 4112
rect -1360 3697 -1199 3768
rect -1128 3697 -1015 3768
rect -1360 3398 -1015 3697
rect -1360 3327 -1195 3398
rect -1124 3327 -1015 3398
rect -1360 3047 -1015 3327
rect -1237 3046 -1015 3047
rect -915 7777 -570 7837
rect -915 7706 -756 7777
rect -685 7706 -570 7777
rect -915 7458 -570 7706
rect -915 7387 -752 7458
rect -681 7387 -570 7458
rect -915 7132 -570 7387
rect -915 7061 -749 7132
rect -678 7061 -570 7132
rect -915 6881 -570 7061
rect -915 6810 -752 6881
rect -681 6810 -570 6881
rect -915 6603 -570 6810
rect -915 6532 -752 6603
rect -681 6532 -570 6603
rect -915 6352 -570 6532
rect -915 6281 -752 6352
rect -681 6281 -570 6352
rect -915 6030 -570 6281
rect -915 5959 -756 6030
rect -685 5959 -570 6030
rect -915 5689 -570 5959
rect -915 5618 -749 5689
rect -678 5618 -570 5689
rect -915 5306 -570 5618
rect -915 5235 -754 5306
rect -683 5235 -570 5306
rect -915 4944 -570 5235
rect -915 4873 -754 4944
rect -683 4873 -570 4944
rect -915 4601 -570 4873
rect -915 4530 -747 4601
rect -676 4530 -570 4601
rect -915 4183 -570 4530
rect -915 4112 -758 4183
rect -687 4112 -570 4183
rect -915 3768 -570 4112
rect -915 3697 -754 3768
rect -683 3697 -570 3768
rect -915 3398 -570 3697
rect -915 3327 -750 3398
rect -679 3327 -570 3398
rect -915 3046 -570 3327
rect -470 7777 -125 7837
rect -470 7706 -311 7777
rect -240 7706 -125 7777
rect -470 7458 -125 7706
rect -470 7387 -307 7458
rect -236 7387 -125 7458
rect -470 7132 -125 7387
rect -470 7061 -304 7132
rect -233 7061 -125 7132
rect -470 6881 -125 7061
rect -470 6810 -307 6881
rect -236 6810 -125 6881
rect -470 6603 -125 6810
rect -470 6532 -307 6603
rect -236 6532 -125 6603
rect -470 6352 -125 6532
rect -470 6281 -307 6352
rect -236 6281 -125 6352
rect -470 6030 -125 6281
rect -470 5959 -311 6030
rect -240 5959 -125 6030
rect -470 5689 -125 5959
rect -470 5618 -304 5689
rect -233 5618 -125 5689
rect -470 5306 -125 5618
rect -470 5235 -309 5306
rect -238 5235 -125 5306
rect -470 4944 -125 5235
rect -470 4873 -309 4944
rect -238 4873 -125 4944
rect -470 4601 -125 4873
rect -470 4530 -302 4601
rect -231 4530 -125 4601
rect -470 4183 -125 4530
rect -470 4112 -313 4183
rect -242 4112 -125 4183
rect -470 3768 -125 4112
rect -470 3697 -309 3768
rect -238 3697 -125 3768
rect -470 3398 -125 3697
rect -470 3327 -305 3398
rect -234 3327 -125 3398
rect -470 3046 -125 3327
rect -25 7777 320 7837
rect -25 7706 134 7777
rect 205 7706 320 7777
rect -25 7458 320 7706
rect -25 7387 138 7458
rect 209 7387 320 7458
rect -25 7132 320 7387
rect -25 7061 141 7132
rect 212 7061 320 7132
rect -25 6881 320 7061
rect -25 6810 138 6881
rect 209 6810 320 6881
rect -25 6603 320 6810
rect -25 6532 138 6603
rect 209 6532 320 6603
rect -25 6352 320 6532
rect -25 6281 138 6352
rect 209 6281 320 6352
rect -25 6030 320 6281
rect -25 5959 134 6030
rect 205 5959 320 6030
rect -25 5689 320 5959
rect -25 5618 141 5689
rect 212 5618 320 5689
rect -25 5306 320 5618
rect -25 5235 136 5306
rect 207 5235 320 5306
rect -25 4944 320 5235
rect -25 4873 136 4944
rect 207 4873 320 4944
rect -25 4601 320 4873
rect -25 4530 143 4601
rect 214 4530 320 4601
rect -25 4183 320 4530
rect -25 4112 132 4183
rect 203 4112 320 4183
rect -25 3768 320 4112
rect -25 3697 136 3768
rect 207 3697 320 3768
rect -25 3398 320 3697
rect -25 3327 140 3398
rect 211 3327 320 3398
rect -25 3046 320 3327
rect 420 7777 765 7837
rect 420 7706 579 7777
rect 650 7706 765 7777
rect 420 7458 765 7706
rect 420 7387 583 7458
rect 654 7387 765 7458
rect 420 7132 765 7387
rect 420 7061 586 7132
rect 657 7061 765 7132
rect 420 6881 765 7061
rect 420 6810 583 6881
rect 654 6810 765 6881
rect 420 6603 765 6810
rect 420 6532 583 6603
rect 654 6532 765 6603
rect 420 6352 765 6532
rect 420 6281 583 6352
rect 654 6281 765 6352
rect 420 6030 765 6281
rect 420 5959 579 6030
rect 650 5959 765 6030
rect 420 5689 765 5959
rect 420 5618 586 5689
rect 657 5618 765 5689
rect 420 5306 765 5618
rect 420 5235 581 5306
rect 652 5235 765 5306
rect 420 4944 765 5235
rect 420 4873 581 4944
rect 652 4873 765 4944
rect 420 4601 765 4873
rect 420 4530 588 4601
rect 659 4530 765 4601
rect 420 4183 765 4530
rect 420 4112 577 4183
rect 648 4112 765 4183
rect 420 3768 765 4112
rect 420 3697 581 3768
rect 652 3697 765 3768
rect 420 3398 765 3697
rect 420 3327 585 3398
rect 656 3327 765 3398
rect 420 3046 765 3327
rect 865 7777 1210 7837
rect 865 7706 1024 7777
rect 1095 7706 1210 7777
rect 865 7458 1210 7706
rect 865 7387 1028 7458
rect 1099 7387 1210 7458
rect 865 7132 1210 7387
rect 865 7061 1031 7132
rect 1102 7061 1210 7132
rect 865 6881 1210 7061
rect 865 6810 1028 6881
rect 1099 6810 1210 6881
rect 865 6603 1210 6810
rect 865 6532 1028 6603
rect 1099 6532 1210 6603
rect 865 6352 1210 6532
rect 865 6281 1028 6352
rect 1099 6281 1210 6352
rect 865 6030 1210 6281
rect 865 5959 1024 6030
rect 1095 5959 1210 6030
rect 865 5689 1210 5959
rect 865 5618 1031 5689
rect 1102 5618 1210 5689
rect 865 5306 1210 5618
rect 865 5235 1026 5306
rect 1097 5235 1210 5306
rect 865 4944 1210 5235
rect 865 4873 1026 4944
rect 1097 4873 1210 4944
rect 865 4601 1210 4873
rect 865 4530 1033 4601
rect 1104 4530 1210 4601
rect 865 4183 1210 4530
rect 865 4112 1022 4183
rect 1093 4112 1210 4183
rect 865 3768 1210 4112
rect 865 3697 1026 3768
rect 1097 3697 1210 3768
rect 865 3398 1210 3697
rect 865 3327 1030 3398
rect 1101 3327 1210 3398
rect 865 3046 1210 3327
rect 1310 7777 1655 7837
rect 1310 7706 1469 7777
rect 1540 7706 1655 7777
rect 1310 7458 1655 7706
rect 1310 7387 1473 7458
rect 1544 7387 1655 7458
rect 1310 7132 1655 7387
rect 1310 7061 1476 7132
rect 1547 7061 1655 7132
rect 1310 6881 1655 7061
rect 1310 6810 1473 6881
rect 1544 6810 1655 6881
rect 1310 6603 1655 6810
rect 1310 6532 1473 6603
rect 1544 6532 1655 6603
rect 1310 6352 1655 6532
rect 1310 6281 1473 6352
rect 1544 6281 1655 6352
rect 1310 6030 1655 6281
rect 1310 5959 1469 6030
rect 1540 5959 1655 6030
rect 1310 5689 1655 5959
rect 1310 5618 1476 5689
rect 1547 5618 1655 5689
rect 1310 5306 1655 5618
rect 1310 5235 1471 5306
rect 1542 5235 1655 5306
rect 1310 4944 1655 5235
rect 1310 4873 1471 4944
rect 1542 4873 1655 4944
rect 1310 4601 1655 4873
rect 1310 4530 1478 4601
rect 1549 4530 1655 4601
rect 1310 4183 1655 4530
rect 1310 4112 1467 4183
rect 1538 4112 1655 4183
rect 1310 3768 1655 4112
rect 1310 3697 1471 3768
rect 1542 3697 1655 3768
rect 1310 3398 1655 3697
rect 1310 3327 1475 3398
rect 1546 3327 1655 3398
rect 1310 3046 1655 3327
rect 1755 7777 2100 7837
rect 1755 7706 1914 7777
rect 1985 7706 2100 7777
rect 1755 7458 2100 7706
rect 1755 7387 1918 7458
rect 1989 7387 2100 7458
rect 1755 7132 2100 7387
rect 1755 7061 1921 7132
rect 1992 7061 2100 7132
rect 1755 6881 2100 7061
rect 1755 6810 1918 6881
rect 1989 6810 2100 6881
rect 1755 6603 2100 6810
rect 1755 6532 1918 6603
rect 1989 6532 2100 6603
rect 1755 6352 2100 6532
rect 1755 6281 1918 6352
rect 1989 6281 2100 6352
rect 1755 6030 2100 6281
rect 1755 5959 1914 6030
rect 1985 5959 2100 6030
rect 1755 5689 2100 5959
rect 1755 5618 1921 5689
rect 1992 5618 2100 5689
rect 1755 5306 2100 5618
rect 1755 5235 1916 5306
rect 1987 5235 2100 5306
rect 1755 4944 2100 5235
rect 1755 4873 1916 4944
rect 1987 4873 2100 4944
rect 1755 4601 2100 4873
rect 1755 4530 1923 4601
rect 1994 4530 2100 4601
rect 1755 4183 2100 4530
rect 1755 4112 1912 4183
rect 1983 4112 2100 4183
rect 1755 3768 2100 4112
rect 1755 3697 1916 3768
rect 1987 3697 2100 3768
rect 1755 3398 2100 3697
rect 1755 3327 1920 3398
rect 1991 3327 2100 3398
rect 1755 3046 2100 3327
rect 2200 7777 2545 7837
rect 2200 7706 2359 7777
rect 2430 7706 2545 7777
rect 2200 7458 2545 7706
rect 2200 7387 2363 7458
rect 2434 7387 2545 7458
rect 2200 7132 2545 7387
rect 2200 7061 2366 7132
rect 2437 7061 2545 7132
rect 2200 6881 2545 7061
rect 2200 6810 2363 6881
rect 2434 6810 2545 6881
rect 2200 6603 2545 6810
rect 2200 6532 2363 6603
rect 2434 6532 2545 6603
rect 2200 6352 2545 6532
rect 2200 6281 2363 6352
rect 2434 6281 2545 6352
rect 2200 6030 2545 6281
rect 2200 5959 2359 6030
rect 2430 5959 2545 6030
rect 2200 5689 2545 5959
rect 2200 5618 2366 5689
rect 2437 5618 2545 5689
rect 2200 5306 2545 5618
rect 2200 5235 2361 5306
rect 2432 5235 2545 5306
rect 2200 4944 2545 5235
rect 2200 4873 2361 4944
rect 2432 4873 2545 4944
rect 2200 4601 2545 4873
rect 2200 4530 2368 4601
rect 2439 4530 2545 4601
rect 2200 4183 2545 4530
rect 2200 4112 2357 4183
rect 2428 4112 2545 4183
rect 2200 3768 2545 4112
rect 2200 3697 2361 3768
rect 2432 3697 2545 3768
rect 2200 3398 2545 3697
rect 2200 3327 2365 3398
rect 2436 3327 2545 3398
rect 2200 3046 2545 3327
rect 2645 7777 3098 7837
rect 2645 7706 2804 7777
rect 2875 7706 3098 7777
rect 2645 7458 3098 7706
rect 2645 7387 2808 7458
rect 2879 7387 3098 7458
rect 2645 7132 3098 7387
rect 2645 7061 2811 7132
rect 2882 7061 3098 7132
rect 2645 6881 3098 7061
rect 2645 6810 2808 6881
rect 2879 6810 3098 6881
rect 2645 6603 3098 6810
rect 2645 6532 2808 6603
rect 2879 6532 3098 6603
rect 2645 6352 3098 6532
rect 2645 6281 2808 6352
rect 2879 6281 3098 6352
rect 2645 6030 3098 6281
rect 2645 5959 2804 6030
rect 2875 5959 3098 6030
rect 2645 5689 3098 5959
rect 2645 5618 2811 5689
rect 2882 5618 3098 5689
rect 2645 5306 3098 5618
rect 2645 5235 2806 5306
rect 2877 5235 3098 5306
rect 2645 4944 3098 5235
rect 2645 4873 2806 4944
rect 2877 4873 3098 4944
rect 2645 4601 3098 4873
rect 2645 4530 2813 4601
rect 2884 4530 3098 4601
rect 2645 4183 3098 4530
rect 2645 4112 2802 4183
rect 2873 4112 3098 4183
rect 2645 3768 3098 4112
rect 2645 3697 2806 3768
rect 2877 3697 3098 3768
rect 2645 3398 3098 3697
rect 2645 3327 2810 3398
rect 2881 3327 3098 3398
rect 2645 3062 3098 3327
rect 2645 3046 3099 3062
<< ndiffc >>
rect -232 506 -132 606
rect -234 273 -134 373
rect 228 506 328 606
rect 226 273 326 373
rect 668 508 768 608
rect 666 275 766 375
rect 1132 508 1232 608
rect 1130 275 1230 375
rect 1558 510 1658 610
rect 1556 277 1656 377
rect 1953 510 2053 610
rect 1951 277 2051 377
<< pdiffc >>
rect -7628 7707 -7557 7778
rect -7624 7388 -7553 7459
rect -7621 7062 -7550 7133
rect -7624 6811 -7553 6882
rect -7624 6533 -7553 6604
rect -7624 6282 -7553 6353
rect -7628 5960 -7557 6031
rect -7621 5619 -7550 5690
rect -7626 5236 -7555 5307
rect -7626 4874 -7555 4945
rect -7619 4531 -7548 4602
rect -7630 4113 -7559 4184
rect -7626 3698 -7555 3769
rect -7622 3328 -7551 3399
rect -7201 7706 -7130 7777
rect -7197 7387 -7126 7458
rect -7194 7061 -7123 7132
rect -7197 6810 -7126 6881
rect -7197 6532 -7126 6603
rect -7197 6281 -7126 6352
rect -7201 5959 -7130 6030
rect -7194 5618 -7123 5689
rect -7199 5235 -7128 5306
rect -7199 4873 -7128 4944
rect -7192 4530 -7121 4601
rect -7203 4112 -7132 4183
rect -7199 3697 -7128 3768
rect -7195 3327 -7124 3398
rect -6756 7706 -6685 7777
rect -6752 7387 -6681 7458
rect -6749 7061 -6678 7132
rect -6752 6810 -6681 6881
rect -6752 6532 -6681 6603
rect -6752 6281 -6681 6352
rect -6756 5959 -6685 6030
rect -6749 5618 -6678 5689
rect -6754 5235 -6683 5306
rect -6754 4873 -6683 4944
rect -6747 4530 -6676 4601
rect -6758 4112 -6687 4183
rect -6754 3697 -6683 3768
rect -6750 3327 -6679 3398
rect -6311 7706 -6240 7777
rect -6307 7387 -6236 7458
rect -6304 7061 -6233 7132
rect -6307 6810 -6236 6881
rect -6307 6532 -6236 6603
rect -6307 6281 -6236 6352
rect -6311 5959 -6240 6030
rect -6304 5618 -6233 5689
rect -6309 5235 -6238 5306
rect -6309 4873 -6238 4944
rect -6302 4530 -6231 4601
rect -6313 4112 -6242 4183
rect -6309 3697 -6238 3768
rect -6305 3327 -6234 3398
rect -5866 7706 -5795 7777
rect -5862 7387 -5791 7458
rect -5859 7061 -5788 7132
rect -5862 6810 -5791 6881
rect -5862 6532 -5791 6603
rect -5862 6281 -5791 6352
rect -5866 5959 -5795 6030
rect -5859 5618 -5788 5689
rect -5864 5235 -5793 5306
rect -5864 4873 -5793 4944
rect -5857 4530 -5786 4601
rect -5868 4112 -5797 4183
rect -5864 3697 -5793 3768
rect -5860 3327 -5789 3398
rect -5421 7706 -5350 7777
rect -5417 7387 -5346 7458
rect -5414 7061 -5343 7132
rect -5417 6810 -5346 6881
rect -5417 6532 -5346 6603
rect -5417 6281 -5346 6352
rect -5421 5959 -5350 6030
rect -5414 5618 -5343 5689
rect -5419 5235 -5348 5306
rect -5419 4873 -5348 4944
rect -5412 4530 -5341 4601
rect -5423 4112 -5352 4183
rect -5419 3697 -5348 3768
rect -5415 3327 -5344 3398
rect -4976 7706 -4905 7777
rect -4972 7387 -4901 7458
rect -4969 7061 -4898 7132
rect -4972 6810 -4901 6881
rect -4972 6532 -4901 6603
rect -4972 6281 -4901 6352
rect -4976 5959 -4905 6030
rect -4969 5618 -4898 5689
rect -4974 5235 -4903 5306
rect -4974 4873 -4903 4944
rect -4967 4530 -4896 4601
rect -4978 4112 -4907 4183
rect -4974 3697 -4903 3768
rect -4970 3327 -4899 3398
rect -4531 7706 -4460 7777
rect -4527 7387 -4456 7458
rect -4524 7061 -4453 7132
rect -4527 6810 -4456 6881
rect -4527 6532 -4456 6603
rect -4527 6281 -4456 6352
rect -4531 5959 -4460 6030
rect -4524 5618 -4453 5689
rect -4529 5235 -4458 5306
rect -4529 4873 -4458 4944
rect -4522 4530 -4451 4601
rect -4533 4112 -4462 4183
rect -4529 3697 -4458 3768
rect -4525 3327 -4454 3398
rect -4086 7706 -4015 7777
rect -4082 7387 -4011 7458
rect -4079 7061 -4008 7132
rect -4082 6810 -4011 6881
rect -4082 6532 -4011 6603
rect -4082 6281 -4011 6352
rect -4086 5959 -4015 6030
rect -4079 5618 -4008 5689
rect -4084 5235 -4013 5306
rect -4084 4873 -4013 4944
rect -4077 4530 -4006 4601
rect -4088 4112 -4017 4183
rect -4084 3697 -4013 3768
rect -4080 3327 -4009 3398
rect -3641 7706 -3570 7777
rect -3637 7387 -3566 7458
rect -3634 7061 -3563 7132
rect -3637 6810 -3566 6881
rect -3637 6532 -3566 6603
rect -3637 6281 -3566 6352
rect -3641 5959 -3570 6030
rect -3634 5618 -3563 5689
rect -3639 5235 -3568 5306
rect -3639 4873 -3568 4944
rect -3632 4530 -3561 4601
rect -3643 4112 -3572 4183
rect -3639 3697 -3568 3768
rect -3635 3327 -3564 3398
rect -3196 7706 -3125 7777
rect -3192 7387 -3121 7458
rect -3189 7061 -3118 7132
rect -3192 6810 -3121 6881
rect -3192 6532 -3121 6603
rect -3192 6281 -3121 6352
rect -3196 5959 -3125 6030
rect -3189 5618 -3118 5689
rect -3194 5235 -3123 5306
rect -3194 4873 -3123 4944
rect -3187 4530 -3116 4601
rect -3198 4112 -3127 4183
rect -3194 3697 -3123 3768
rect -3190 3327 -3119 3398
rect -1628 7707 -1557 7778
rect -1624 7388 -1553 7459
rect -1621 7062 -1550 7133
rect -1624 6811 -1553 6882
rect -1624 6533 -1553 6604
rect -1624 6282 -1553 6353
rect -1628 5960 -1557 6031
rect -1621 5619 -1550 5690
rect -1626 5236 -1555 5307
rect -1626 4874 -1555 4945
rect -1619 4531 -1548 4602
rect -1630 4113 -1559 4184
rect -1626 3698 -1555 3769
rect -1622 3328 -1551 3399
rect -1201 7706 -1130 7777
rect -1197 7387 -1126 7458
rect -1194 7061 -1123 7132
rect -1197 6810 -1126 6881
rect -1197 6532 -1126 6603
rect -1197 6281 -1126 6352
rect -1201 5959 -1130 6030
rect -1194 5618 -1123 5689
rect -1199 5235 -1128 5306
rect -1199 4873 -1128 4944
rect -1192 4530 -1121 4601
rect -1203 4112 -1132 4183
rect -1199 3697 -1128 3768
rect -1195 3327 -1124 3398
rect -756 7706 -685 7777
rect -752 7387 -681 7458
rect -749 7061 -678 7132
rect -752 6810 -681 6881
rect -752 6532 -681 6603
rect -752 6281 -681 6352
rect -756 5959 -685 6030
rect -749 5618 -678 5689
rect -754 5235 -683 5306
rect -754 4873 -683 4944
rect -747 4530 -676 4601
rect -758 4112 -687 4183
rect -754 3697 -683 3768
rect -750 3327 -679 3398
rect -311 7706 -240 7777
rect -307 7387 -236 7458
rect -304 7061 -233 7132
rect -307 6810 -236 6881
rect -307 6532 -236 6603
rect -307 6281 -236 6352
rect -311 5959 -240 6030
rect -304 5618 -233 5689
rect -309 5235 -238 5306
rect -309 4873 -238 4944
rect -302 4530 -231 4601
rect -313 4112 -242 4183
rect -309 3697 -238 3768
rect -305 3327 -234 3398
rect 134 7706 205 7777
rect 138 7387 209 7458
rect 141 7061 212 7132
rect 138 6810 209 6881
rect 138 6532 209 6603
rect 138 6281 209 6352
rect 134 5959 205 6030
rect 141 5618 212 5689
rect 136 5235 207 5306
rect 136 4873 207 4944
rect 143 4530 214 4601
rect 132 4112 203 4183
rect 136 3697 207 3768
rect 140 3327 211 3398
rect 579 7706 650 7777
rect 583 7387 654 7458
rect 586 7061 657 7132
rect 583 6810 654 6881
rect 583 6532 654 6603
rect 583 6281 654 6352
rect 579 5959 650 6030
rect 586 5618 657 5689
rect 581 5235 652 5306
rect 581 4873 652 4944
rect 588 4530 659 4601
rect 577 4112 648 4183
rect 581 3697 652 3768
rect 585 3327 656 3398
rect 1024 7706 1095 7777
rect 1028 7387 1099 7458
rect 1031 7061 1102 7132
rect 1028 6810 1099 6881
rect 1028 6532 1099 6603
rect 1028 6281 1099 6352
rect 1024 5959 1095 6030
rect 1031 5618 1102 5689
rect 1026 5235 1097 5306
rect 1026 4873 1097 4944
rect 1033 4530 1104 4601
rect 1022 4112 1093 4183
rect 1026 3697 1097 3768
rect 1030 3327 1101 3398
rect 1469 7706 1540 7777
rect 1473 7387 1544 7458
rect 1476 7061 1547 7132
rect 1473 6810 1544 6881
rect 1473 6532 1544 6603
rect 1473 6281 1544 6352
rect 1469 5959 1540 6030
rect 1476 5618 1547 5689
rect 1471 5235 1542 5306
rect 1471 4873 1542 4944
rect 1478 4530 1549 4601
rect 1467 4112 1538 4183
rect 1471 3697 1542 3768
rect 1475 3327 1546 3398
rect 1914 7706 1985 7777
rect 1918 7387 1989 7458
rect 1921 7061 1992 7132
rect 1918 6810 1989 6881
rect 1918 6532 1989 6603
rect 1918 6281 1989 6352
rect 1914 5959 1985 6030
rect 1921 5618 1992 5689
rect 1916 5235 1987 5306
rect 1916 4873 1987 4944
rect 1923 4530 1994 4601
rect 1912 4112 1983 4183
rect 1916 3697 1987 3768
rect 1920 3327 1991 3398
rect 2359 7706 2430 7777
rect 2363 7387 2434 7458
rect 2366 7061 2437 7132
rect 2363 6810 2434 6881
rect 2363 6532 2434 6603
rect 2363 6281 2434 6352
rect 2359 5959 2430 6030
rect 2366 5618 2437 5689
rect 2361 5235 2432 5306
rect 2361 4873 2432 4944
rect 2368 4530 2439 4601
rect 2357 4112 2428 4183
rect 2361 3697 2432 3768
rect 2365 3327 2436 3398
rect 2804 7706 2875 7777
rect 2808 7387 2879 7458
rect 2811 7061 2882 7132
rect 2808 6810 2879 6881
rect 2808 6532 2879 6603
rect 2808 6281 2879 6352
rect 2804 5959 2875 6030
rect 2811 5618 2882 5689
rect 2806 5235 2877 5306
rect 2806 4873 2877 4944
rect 2813 4530 2884 4601
rect 2802 4112 2873 4183
rect 2806 3697 2877 3768
rect 2810 3327 2881 3398
<< poly >>
rect -7460 7837 -7360 8159
rect -7015 7837 -6915 8159
rect -6570 7837 -6470 8159
rect -6125 7837 -6025 8159
rect -5680 7837 -5580 8159
rect -5235 7837 -5135 8159
rect -4790 7837 -4690 8159
rect -4345 7837 -4245 8159
rect -3900 7837 -3800 8159
rect -3455 7837 -3355 8159
rect -1460 7837 -1360 8159
rect -1015 7837 -915 8159
rect -570 7837 -470 8159
rect -125 7837 -25 8159
rect 320 7837 420 8159
rect 765 7837 865 8159
rect 1210 7837 1310 8159
rect 1655 7837 1755 8159
rect 2100 7837 2200 8159
rect 2545 7837 2645 8159
rect -7460 2755 -7360 3047
rect -7015 2755 -6915 3046
rect -6570 2755 -6470 3046
rect -6125 2755 -6025 3046
rect -5680 2755 -5580 3046
rect -5235 2755 -5135 3046
rect -4790 2755 -4690 3046
rect -4345 2755 -4245 3046
rect -3900 2755 -3800 3046
rect -3455 2755 -3355 3046
rect -7460 2753 -2908 2755
rect -2473 2753 -2112 2768
rect -1460 2753 -1360 3047
rect -1015 2753 -915 3046
rect -570 2753 -470 3046
rect -125 2753 -25 3046
rect 320 2753 420 3046
rect 765 2753 865 3046
rect 1210 2753 1310 3046
rect 1655 2753 1755 3046
rect 2100 2753 2200 3046
rect 2545 2753 2645 3046
rect -7460 2655 -2461 2753
rect -7013 2653 -2461 2655
rect -2473 2406 -2461 2653
rect -2131 2655 2645 2753
rect -2131 2653 2200 2655
rect -2131 2406 -2112 2653
rect -2473 2396 -2112 2406
rect -1003 1185 -603 1193
rect -1003 813 -986 1185
rect -625 1045 -603 1185
rect -625 1043 1115 1045
rect -625 945 1848 1043
rect -625 813 -603 945
rect 0 943 1848 945
rect 0 847 100 943
rect 457 847 557 943
rect 905 847 1005 943
rect 1353 847 1453 943
rect 1746 847 1846 943
rect -1003 793 -603 813
rect 0 -196 100 -13
rect 457 -196 557 -13
rect 905 -196 1005 -13
rect 1353 -205 1453 -13
rect 1746 -196 1846 -13
<< polycont >>
rect -2461 2406 -2131 2753
rect -986 813 -625 1185
<< locali >>
rect -7210 8717 -3549 8727
rect 309 8726 1068 8727
rect 1827 8726 2452 8727
rect -7210 8714 -3729 8717
rect -7210 8711 -5473 8714
rect -7210 8541 -7194 8711
rect -7024 8708 -5473 8711
rect -7024 8541 -6351 8708
rect -7210 8538 -6351 8541
rect -6181 8544 -5473 8708
rect -5303 8708 -3729 8714
rect -5303 8544 -4578 8708
rect -6181 8538 -4578 8544
rect -4408 8547 -3729 8708
rect -3559 8586 -3549 8717
rect -1208 8716 2452 8726
rect -1208 8706 538 8716
rect -1208 8705 -358 8706
rect -1208 8630 -1198 8705
rect -3559 8547 -3548 8586
rect -4408 8538 -3548 8547
rect -7210 8532 -3548 8538
rect -7210 8530 -5892 8532
rect -5760 8530 -5001 8532
rect -4869 8530 -4110 8532
rect -3978 8530 -3548 8532
rect -7637 7778 -7537 7851
rect -7637 7707 -7628 7778
rect -7557 7707 -7537 7778
rect -7637 7459 -7537 7707
rect -7637 7388 -7624 7459
rect -7553 7388 -7537 7459
rect -7637 7133 -7537 7388
rect -7637 7062 -7621 7133
rect -7550 7062 -7537 7133
rect -7637 6882 -7537 7062
rect -7637 6811 -7624 6882
rect -7553 6811 -7537 6882
rect -7637 6604 -7537 6811
rect -7637 6533 -7624 6604
rect -7553 6533 -7537 6604
rect -7637 6353 -7537 6533
rect -7637 6282 -7624 6353
rect -7553 6282 -7537 6353
rect -7637 6031 -7537 6282
rect -7637 5960 -7628 6031
rect -7557 5960 -7537 6031
rect -7637 5690 -7537 5960
rect -7637 5619 -7621 5690
rect -7550 5619 -7537 5690
rect -7637 5307 -7537 5619
rect -7637 5236 -7626 5307
rect -7555 5236 -7537 5307
rect -7637 4945 -7537 5236
rect -7637 4874 -7626 4945
rect -7555 4874 -7537 4945
rect -7637 4602 -7537 4874
rect -7637 4531 -7619 4602
rect -7548 4531 -7537 4602
rect -7637 4184 -7537 4531
rect -7637 4113 -7630 4184
rect -7559 4113 -7537 4184
rect -7637 3769 -7537 4113
rect -7637 3698 -7626 3769
rect -7555 3698 -7537 3769
rect -7637 3399 -7537 3698
rect -7637 3328 -7622 3399
rect -7551 3328 -7537 3399
rect -7637 2521 -7537 3328
rect -7210 7777 -7110 8530
rect -7210 7706 -7201 7777
rect -7130 7706 -7110 7777
rect -7210 7458 -7110 7706
rect -7210 7387 -7197 7458
rect -7126 7387 -7110 7458
rect -7210 7132 -7110 7387
rect -7210 7061 -7194 7132
rect -7123 7061 -7110 7132
rect -7210 6881 -7110 7061
rect -7210 6810 -7197 6881
rect -7126 6810 -7110 6881
rect -7210 6603 -7110 6810
rect -7210 6532 -7197 6603
rect -7126 6532 -7110 6603
rect -7210 6352 -7110 6532
rect -7210 6281 -7197 6352
rect -7126 6281 -7110 6352
rect -7210 6030 -7110 6281
rect -7210 5959 -7201 6030
rect -7130 5959 -7110 6030
rect -7210 5689 -7110 5959
rect -7210 5618 -7194 5689
rect -7123 5618 -7110 5689
rect -7210 5306 -7110 5618
rect -7210 5235 -7199 5306
rect -7128 5235 -7110 5306
rect -7210 4944 -7110 5235
rect -7210 4873 -7199 4944
rect -7128 4873 -7110 4944
rect -7210 4601 -7110 4873
rect -7210 4530 -7192 4601
rect -7121 4530 -7110 4601
rect -7210 4183 -7110 4530
rect -7210 4112 -7203 4183
rect -7132 4112 -7110 4183
rect -7210 3768 -7110 4112
rect -7210 3697 -7199 3768
rect -7128 3697 -7110 3768
rect -7210 3398 -7110 3697
rect -7210 3327 -7195 3398
rect -7124 3327 -7110 3398
rect -7210 3060 -7110 3327
rect -6765 7777 -6665 7837
rect -6765 7706 -6756 7777
rect -6685 7706 -6665 7777
rect -6765 7458 -6665 7706
rect -6765 7387 -6752 7458
rect -6681 7387 -6665 7458
rect -6765 7132 -6665 7387
rect -6765 7061 -6749 7132
rect -6678 7061 -6665 7132
rect -6765 6881 -6665 7061
rect -6765 6810 -6752 6881
rect -6681 6810 -6665 6881
rect -6765 6603 -6665 6810
rect -6765 6532 -6752 6603
rect -6681 6532 -6665 6603
rect -6765 6352 -6665 6532
rect -6765 6281 -6752 6352
rect -6681 6281 -6665 6352
rect -6765 6030 -6665 6281
rect -6765 5959 -6756 6030
rect -6685 5959 -6665 6030
rect -6765 5689 -6665 5959
rect -6765 5618 -6749 5689
rect -6678 5618 -6665 5689
rect -6765 5306 -6665 5618
rect -6765 5235 -6754 5306
rect -6683 5235 -6665 5306
rect -6765 4944 -6665 5235
rect -6765 4873 -6754 4944
rect -6683 4873 -6665 4944
rect -6765 4601 -6665 4873
rect -6765 4530 -6747 4601
rect -6676 4530 -6665 4601
rect -6765 4183 -6665 4530
rect -6765 4112 -6758 4183
rect -6687 4112 -6665 4183
rect -6765 3768 -6665 4112
rect -6765 3697 -6754 3768
rect -6683 3697 -6665 3768
rect -6765 3398 -6665 3697
rect -6765 3327 -6750 3398
rect -6679 3328 -6665 3398
rect -6320 7777 -6220 8530
rect -6320 7706 -6311 7777
rect -6240 7706 -6220 7777
rect -6320 7458 -6220 7706
rect -6320 7387 -6307 7458
rect -6236 7387 -6220 7458
rect -6320 7132 -6220 7387
rect -6320 7061 -6304 7132
rect -6233 7061 -6220 7132
rect -6320 6881 -6220 7061
rect -6320 6810 -6307 6881
rect -6236 6810 -6220 6881
rect -6320 6603 -6220 6810
rect -6320 6532 -6307 6603
rect -6236 6532 -6220 6603
rect -6320 6352 -6220 6532
rect -6320 6281 -6307 6352
rect -6236 6281 -6220 6352
rect -6320 6030 -6220 6281
rect -6320 5959 -6311 6030
rect -6240 5959 -6220 6030
rect -6320 5689 -6220 5959
rect -6320 5618 -6304 5689
rect -6233 5618 -6220 5689
rect -6320 5306 -6220 5618
rect -6320 5235 -6309 5306
rect -6238 5235 -6220 5306
rect -6320 4944 -6220 5235
rect -6320 4873 -6309 4944
rect -6238 4873 -6220 4944
rect -6320 4601 -6220 4873
rect -6320 4530 -6302 4601
rect -6231 4530 -6220 4601
rect -6320 4183 -6220 4530
rect -6320 4112 -6313 4183
rect -6242 4112 -6220 4183
rect -6320 3768 -6220 4112
rect -6320 3697 -6309 3768
rect -6238 3697 -6220 3768
rect -6320 3398 -6220 3697
rect -6679 3327 -6664 3328
rect -6765 3060 -6664 3327
rect -6320 3327 -6305 3398
rect -6234 3327 -6220 3398
rect -6320 3060 -6220 3327
rect -5875 7777 -5775 7833
rect -5875 7706 -5866 7777
rect -5795 7706 -5775 7777
rect -5875 7458 -5775 7706
rect -5875 7387 -5862 7458
rect -5791 7387 -5775 7458
rect -5875 7132 -5775 7387
rect -5875 7061 -5859 7132
rect -5788 7061 -5775 7132
rect -5875 6881 -5775 7061
rect -5875 6810 -5862 6881
rect -5791 6810 -5775 6881
rect -5875 6603 -5775 6810
rect -5875 6532 -5862 6603
rect -5791 6532 -5775 6603
rect -5875 6352 -5775 6532
rect -5875 6281 -5862 6352
rect -5791 6281 -5775 6352
rect -5875 6030 -5775 6281
rect -5875 5959 -5866 6030
rect -5795 5959 -5775 6030
rect -5875 5689 -5775 5959
rect -5875 5618 -5859 5689
rect -5788 5618 -5775 5689
rect -5875 5306 -5775 5618
rect -5875 5235 -5864 5306
rect -5793 5235 -5775 5306
rect -5875 4944 -5775 5235
rect -5875 4873 -5864 4944
rect -5793 4873 -5775 4944
rect -5875 4601 -5775 4873
rect -5875 4530 -5857 4601
rect -5786 4530 -5775 4601
rect -5875 4183 -5775 4530
rect -5875 4112 -5868 4183
rect -5797 4112 -5775 4183
rect -5875 3768 -5775 4112
rect -5875 3697 -5864 3768
rect -5793 3697 -5775 3768
rect -5875 3398 -5775 3697
rect -5875 3327 -5860 3398
rect -5789 3327 -5775 3398
rect -6764 2521 -6664 3060
rect -5875 2521 -5775 3327
rect -5430 7777 -5330 8530
rect -5430 7706 -5421 7777
rect -5350 7706 -5330 7777
rect -5430 7458 -5330 7706
rect -5430 7387 -5417 7458
rect -5346 7387 -5330 7458
rect -5430 7132 -5330 7387
rect -5430 7061 -5414 7132
rect -5343 7061 -5330 7132
rect -5430 6881 -5330 7061
rect -5430 6810 -5417 6881
rect -5346 6810 -5330 6881
rect -5430 6603 -5330 6810
rect -5430 6532 -5417 6603
rect -5346 6532 -5330 6603
rect -5430 6352 -5330 6532
rect -5430 6281 -5417 6352
rect -5346 6281 -5330 6352
rect -5430 6030 -5330 6281
rect -5430 5959 -5421 6030
rect -5350 5959 -5330 6030
rect -5430 5689 -5330 5959
rect -5430 5618 -5414 5689
rect -5343 5618 -5330 5689
rect -5430 5306 -5330 5618
rect -5430 5235 -5419 5306
rect -5348 5235 -5330 5306
rect -5430 4944 -5330 5235
rect -5430 4873 -5419 4944
rect -5348 4873 -5330 4944
rect -5430 4601 -5330 4873
rect -5430 4530 -5412 4601
rect -5341 4530 -5330 4601
rect -5430 4183 -5330 4530
rect -5430 4112 -5423 4183
rect -5352 4112 -5330 4183
rect -5430 3768 -5330 4112
rect -5430 3697 -5419 3768
rect -5348 3697 -5330 3768
rect -5430 3398 -5330 3697
rect -5430 3327 -5415 3398
rect -5344 3327 -5330 3398
rect -5430 3060 -5330 3327
rect -4985 7777 -4885 7833
rect -4985 7706 -4976 7777
rect -4905 7706 -4885 7777
rect -4985 7458 -4885 7706
rect -4985 7387 -4972 7458
rect -4901 7387 -4885 7458
rect -4985 7132 -4885 7387
rect -4985 7061 -4969 7132
rect -4898 7061 -4885 7132
rect -4985 6881 -4885 7061
rect -4985 6810 -4972 6881
rect -4901 6810 -4885 6881
rect -4985 6603 -4885 6810
rect -4985 6532 -4972 6603
rect -4901 6532 -4885 6603
rect -4985 6352 -4885 6532
rect -4985 6281 -4972 6352
rect -4901 6281 -4885 6352
rect -4985 6030 -4885 6281
rect -4985 5959 -4976 6030
rect -4905 5959 -4885 6030
rect -4985 5689 -4885 5959
rect -4985 5618 -4969 5689
rect -4898 5618 -4885 5689
rect -4985 5306 -4885 5618
rect -4985 5235 -4974 5306
rect -4903 5235 -4885 5306
rect -4985 4944 -4885 5235
rect -4985 4873 -4974 4944
rect -4903 4873 -4885 4944
rect -4985 4601 -4885 4873
rect -4985 4530 -4967 4601
rect -4896 4530 -4885 4601
rect -4985 4183 -4885 4530
rect -4985 4112 -4978 4183
rect -4907 4112 -4885 4183
rect -4985 3768 -4885 4112
rect -4985 3697 -4974 3768
rect -4903 3697 -4885 3768
rect -4985 3398 -4885 3697
rect -4985 3327 -4970 3398
rect -4899 3327 -4885 3398
rect -4540 7777 -4440 8530
rect -3650 8504 -3548 8530
rect -1210 8535 -1198 8630
rect -1028 8536 -358 8705
rect -188 8546 538 8706
rect 708 8713 2452 8716
rect 708 8710 2269 8713
rect 708 8546 1418 8710
rect -188 8540 1418 8546
rect 1588 8543 2269 8710
rect 2439 8543 2452 8713
rect 1588 8540 2452 8543
rect -188 8536 2452 8540
rect -1028 8535 2452 8536
rect -1210 8530 2452 8535
rect -1210 8529 309 8530
rect -4540 7706 -4531 7777
rect -4460 7706 -4440 7777
rect -4540 7458 -4440 7706
rect -4540 7387 -4527 7458
rect -4456 7387 -4440 7458
rect -4540 7132 -4440 7387
rect -4540 7061 -4524 7132
rect -4453 7061 -4440 7132
rect -4540 6881 -4440 7061
rect -4540 6810 -4527 6881
rect -4456 6810 -4440 6881
rect -4540 6603 -4440 6810
rect -4540 6532 -4527 6603
rect -4456 6532 -4440 6603
rect -4540 6352 -4440 6532
rect -4540 6281 -4527 6352
rect -4456 6281 -4440 6352
rect -4540 6030 -4440 6281
rect -4540 5959 -4531 6030
rect -4460 5959 -4440 6030
rect -4540 5689 -4440 5959
rect -4540 5618 -4524 5689
rect -4453 5618 -4440 5689
rect -4540 5306 -4440 5618
rect -4540 5235 -4529 5306
rect -4458 5235 -4440 5306
rect -4540 4944 -4440 5235
rect -4540 4873 -4529 4944
rect -4458 4873 -4440 4944
rect -4540 4601 -4440 4873
rect -4540 4530 -4522 4601
rect -4451 4530 -4440 4601
rect -4540 4183 -4440 4530
rect -4540 4112 -4533 4183
rect -4462 4112 -4440 4183
rect -4540 3768 -4440 4112
rect -4540 3697 -4529 3768
rect -4458 3697 -4440 3768
rect -4540 3398 -4440 3697
rect -4540 3327 -4525 3398
rect -4454 3327 -4440 3398
rect -4985 3060 -4884 3327
rect -4540 3060 -4440 3327
rect -4095 7777 -3995 7833
rect -4095 7706 -4086 7777
rect -4015 7706 -3995 7777
rect -4095 7458 -3995 7706
rect -4095 7387 -4082 7458
rect -4011 7387 -3995 7458
rect -4095 7132 -3995 7387
rect -4095 7061 -4079 7132
rect -4008 7061 -3995 7132
rect -4095 6881 -3995 7061
rect -4095 6810 -4082 6881
rect -4011 6810 -3995 6881
rect -4095 6603 -3995 6810
rect -4095 6532 -4082 6603
rect -4011 6532 -3995 6603
rect -4095 6352 -3995 6532
rect -4095 6281 -4082 6352
rect -4011 6281 -3995 6352
rect -4095 6030 -3995 6281
rect -4095 5959 -4086 6030
rect -4015 5959 -3995 6030
rect -4095 5689 -3995 5959
rect -4095 5618 -4079 5689
rect -4008 5618 -3995 5689
rect -4095 5306 -3995 5618
rect -4095 5235 -4084 5306
rect -4013 5235 -3995 5306
rect -4095 4944 -3995 5235
rect -4095 4873 -4084 4944
rect -4013 4873 -3995 4944
rect -4095 4601 -3995 4873
rect -4095 4530 -4077 4601
rect -4006 4530 -3995 4601
rect -4095 4183 -3995 4530
rect -4095 4112 -4088 4183
rect -4017 4112 -3995 4183
rect -4095 3768 -3995 4112
rect -4095 3697 -4084 3768
rect -4013 3697 -3995 3768
rect -4095 3398 -3995 3697
rect -4095 3327 -4080 3398
rect -4009 3327 -3995 3398
rect -3650 7777 -3550 8504
rect -3650 7706 -3641 7777
rect -3570 7706 -3550 7777
rect -3650 7458 -3550 7706
rect -3650 7387 -3637 7458
rect -3566 7387 -3550 7458
rect -3650 7132 -3550 7387
rect -3650 7061 -3634 7132
rect -3563 7061 -3550 7132
rect -3650 6881 -3550 7061
rect -3650 6810 -3637 6881
rect -3566 6810 -3550 6881
rect -3650 6603 -3550 6810
rect -3650 6532 -3637 6603
rect -3566 6532 -3550 6603
rect -3650 6352 -3550 6532
rect -3650 6281 -3637 6352
rect -3566 6281 -3550 6352
rect -3650 6030 -3550 6281
rect -3650 5959 -3641 6030
rect -3570 5959 -3550 6030
rect -3650 5689 -3550 5959
rect -3650 5618 -3634 5689
rect -3563 5618 -3550 5689
rect -3650 5306 -3550 5618
rect -3650 5235 -3639 5306
rect -3568 5235 -3550 5306
rect -3650 4944 -3550 5235
rect -3650 4873 -3639 4944
rect -3568 4873 -3550 4944
rect -3650 4601 -3550 4873
rect -3650 4530 -3632 4601
rect -3561 4530 -3550 4601
rect -3650 4183 -3550 4530
rect -3650 4112 -3643 4183
rect -3572 4112 -3550 4183
rect -3650 3768 -3550 4112
rect -3650 3697 -3639 3768
rect -3568 3697 -3550 3768
rect -3650 3398 -3550 3697
rect -3650 3327 -3635 3398
rect -3564 3327 -3550 3398
rect -4095 3060 -3993 3327
rect -3650 3060 -3550 3327
rect -3205 7777 -3105 7833
rect -3205 7706 -3196 7777
rect -3125 7706 -3105 7777
rect -3205 7458 -3105 7706
rect -3205 7387 -3192 7458
rect -3121 7387 -3105 7458
rect -3205 7132 -3105 7387
rect -3205 7061 -3189 7132
rect -3118 7061 -3105 7132
rect -3205 6881 -3105 7061
rect -3205 6810 -3192 6881
rect -3121 6810 -3105 6881
rect -3205 6603 -3105 6810
rect -3205 6532 -3192 6603
rect -3121 6532 -3105 6603
rect -3205 6352 -3105 6532
rect -3205 6281 -3192 6352
rect -3121 6281 -3105 6352
rect -3205 6030 -3105 6281
rect -3205 5959 -3196 6030
rect -3125 5959 -3105 6030
rect -3205 5689 -3105 5959
rect -3205 5618 -3189 5689
rect -3118 5618 -3105 5689
rect -3205 5306 -3105 5618
rect -3205 5235 -3194 5306
rect -3123 5235 -3105 5306
rect -3205 4944 -3105 5235
rect -3205 4873 -3194 4944
rect -3123 4873 -3105 4944
rect -3205 4601 -3105 4873
rect -3205 4530 -3187 4601
rect -3116 4530 -3105 4601
rect -3205 4183 -3105 4530
rect -3205 4112 -3198 4183
rect -3127 4112 -3105 4183
rect -3205 3768 -3105 4112
rect -3205 3697 -3194 3768
rect -3123 3697 -3105 3768
rect -3205 3398 -3105 3697
rect -3205 3327 -3190 3398
rect -3119 3327 -3105 3398
rect -1637 7778 -1537 7851
rect -1637 7707 -1628 7778
rect -1557 7707 -1537 7778
rect -1637 7459 -1537 7707
rect -1637 7388 -1624 7459
rect -1553 7388 -1537 7459
rect -1637 7133 -1537 7388
rect -1637 7062 -1621 7133
rect -1550 7062 -1537 7133
rect -1637 6882 -1537 7062
rect -1637 6811 -1624 6882
rect -1553 6811 -1537 6882
rect -1637 6604 -1537 6811
rect -1637 6533 -1624 6604
rect -1553 6533 -1537 6604
rect -1637 6353 -1537 6533
rect -1637 6282 -1624 6353
rect -1553 6282 -1537 6353
rect -1637 6031 -1537 6282
rect -1637 5960 -1628 6031
rect -1557 5960 -1537 6031
rect -1637 5690 -1537 5960
rect -1637 5619 -1621 5690
rect -1550 5619 -1537 5690
rect -1637 5307 -1537 5619
rect -1637 5236 -1626 5307
rect -1555 5236 -1537 5307
rect -1637 4945 -1537 5236
rect -1637 4874 -1626 4945
rect -1555 4874 -1537 4945
rect -1637 4602 -1537 4874
rect -1637 4531 -1619 4602
rect -1548 4531 -1537 4602
rect -1637 4184 -1537 4531
rect -1637 4113 -1630 4184
rect -1559 4113 -1537 4184
rect -1637 3769 -1537 4113
rect -1637 3698 -1626 3769
rect -1555 3698 -1537 3769
rect -1637 3399 -1537 3698
rect -1637 3328 -1622 3399
rect -1551 3328 -1537 3399
rect -3205 3060 -3102 3327
rect -5360 2521 -5228 2524
rect -4984 2521 -4884 3060
rect -4093 2521 -3993 3060
rect -3202 2521 -3102 3060
rect -2473 2753 -2112 2768
rect -2473 2521 -2461 2753
rect -7637 2421 -2461 2521
rect -5360 2409 -5228 2421
rect -2473 2406 -2461 2421
rect -2131 2521 -2112 2753
rect -1637 2521 -1537 3328
rect -1210 7777 -1110 8529
rect -1210 7706 -1201 7777
rect -1130 7706 -1110 7777
rect -1210 7458 -1110 7706
rect -1210 7387 -1197 7458
rect -1126 7387 -1110 7458
rect -1210 7132 -1110 7387
rect -1210 7061 -1194 7132
rect -1123 7061 -1110 7132
rect -1210 6881 -1110 7061
rect -1210 6810 -1197 6881
rect -1126 6810 -1110 6881
rect -1210 6603 -1110 6810
rect -1210 6532 -1197 6603
rect -1126 6532 -1110 6603
rect -1210 6352 -1110 6532
rect -1210 6281 -1197 6352
rect -1126 6281 -1110 6352
rect -1210 6030 -1110 6281
rect -1210 5959 -1201 6030
rect -1130 5959 -1110 6030
rect -1210 5689 -1110 5959
rect -1210 5618 -1194 5689
rect -1123 5618 -1110 5689
rect -1210 5306 -1110 5618
rect -1210 5235 -1199 5306
rect -1128 5235 -1110 5306
rect -1210 4944 -1110 5235
rect -1210 4873 -1199 4944
rect -1128 4873 -1110 4944
rect -1210 4601 -1110 4873
rect -1210 4530 -1192 4601
rect -1121 4530 -1110 4601
rect -1210 4183 -1110 4530
rect -1210 4112 -1203 4183
rect -1132 4112 -1110 4183
rect -1210 3768 -1110 4112
rect -1210 3697 -1199 3768
rect -1128 3697 -1110 3768
rect -1210 3398 -1110 3697
rect -1210 3327 -1195 3398
rect -1124 3327 -1110 3398
rect -1210 3060 -1110 3327
rect -765 7777 -665 7832
rect -765 7706 -756 7777
rect -685 7706 -665 7777
rect -765 7458 -665 7706
rect -765 7387 -752 7458
rect -681 7387 -665 7458
rect -765 7132 -665 7387
rect -765 7061 -749 7132
rect -678 7061 -665 7132
rect -765 6881 -665 7061
rect -765 6810 -752 6881
rect -681 6810 -665 6881
rect -765 6603 -665 6810
rect -765 6532 -752 6603
rect -681 6532 -665 6603
rect -765 6352 -665 6532
rect -765 6281 -752 6352
rect -681 6281 -665 6352
rect -765 6030 -665 6281
rect -765 5959 -756 6030
rect -685 5959 -665 6030
rect -765 5689 -665 5959
rect -765 5618 -749 5689
rect -678 5618 -665 5689
rect -765 5306 -665 5618
rect -765 5235 -754 5306
rect -683 5235 -665 5306
rect -765 4944 -665 5235
rect -765 4873 -754 4944
rect -683 4873 -665 4944
rect -765 4601 -665 4873
rect -765 4530 -747 4601
rect -676 4530 -665 4601
rect -765 4183 -665 4530
rect -765 4112 -758 4183
rect -687 4112 -665 4183
rect -765 3768 -665 4112
rect -765 3697 -754 3768
rect -683 3697 -665 3768
rect -765 3398 -665 3697
rect -765 3327 -750 3398
rect -679 3328 -665 3398
rect -320 7777 -220 8529
rect -320 7706 -311 7777
rect -240 7706 -220 7777
rect -320 7458 -220 7706
rect -320 7387 -307 7458
rect -236 7387 -220 7458
rect -320 7132 -220 7387
rect -320 7061 -304 7132
rect -233 7061 -220 7132
rect -320 6881 -220 7061
rect -320 6810 -307 6881
rect -236 6810 -220 6881
rect -320 6603 -220 6810
rect -320 6532 -307 6603
rect -236 6532 -220 6603
rect -320 6352 -220 6532
rect -320 6281 -307 6352
rect -236 6281 -220 6352
rect -320 6030 -220 6281
rect -320 5959 -311 6030
rect -240 5959 -220 6030
rect -320 5689 -220 5959
rect -320 5618 -304 5689
rect -233 5618 -220 5689
rect -320 5306 -220 5618
rect -320 5235 -309 5306
rect -238 5235 -220 5306
rect -320 4944 -220 5235
rect -320 4873 -309 4944
rect -238 4873 -220 4944
rect -320 4601 -220 4873
rect -320 4530 -302 4601
rect -231 4530 -220 4601
rect -320 4183 -220 4530
rect -320 4112 -313 4183
rect -242 4112 -220 4183
rect -320 3768 -220 4112
rect -320 3697 -309 3768
rect -238 3697 -220 3768
rect -320 3398 -220 3697
rect -679 3327 -664 3328
rect -765 3060 -664 3327
rect -320 3327 -305 3398
rect -234 3327 -220 3398
rect -320 3060 -220 3327
rect 125 7777 225 7833
rect 125 7706 134 7777
rect 205 7706 225 7777
rect 125 7458 225 7706
rect 125 7387 138 7458
rect 209 7387 225 7458
rect 125 7132 225 7387
rect 125 7061 141 7132
rect 212 7061 225 7132
rect 125 6881 225 7061
rect 125 6810 138 6881
rect 209 6810 225 6881
rect 125 6603 225 6810
rect 125 6532 138 6603
rect 209 6532 225 6603
rect 125 6352 225 6532
rect 125 6281 138 6352
rect 209 6281 225 6352
rect 125 6030 225 6281
rect 125 5959 134 6030
rect 205 5959 225 6030
rect 125 5689 225 5959
rect 125 5618 141 5689
rect 212 5618 225 5689
rect 125 5306 225 5618
rect 125 5235 136 5306
rect 207 5235 225 5306
rect 125 4944 225 5235
rect 125 4873 136 4944
rect 207 4873 225 4944
rect 125 4601 225 4873
rect 125 4530 143 4601
rect 214 4530 225 4601
rect 125 4183 225 4530
rect 125 4112 132 4183
rect 203 4112 225 4183
rect 125 3768 225 4112
rect 125 3697 136 3768
rect 207 3697 225 3768
rect 125 3398 225 3697
rect 125 3327 140 3398
rect 211 3327 225 3398
rect -764 2521 -664 3060
rect 125 2521 225 3327
rect 570 7777 670 8530
rect 1068 8529 1827 8530
rect 570 7706 579 7777
rect 650 7706 670 7777
rect 570 7458 670 7706
rect 570 7387 583 7458
rect 654 7387 670 7458
rect 570 7132 670 7387
rect 570 7061 586 7132
rect 657 7061 670 7132
rect 570 6881 670 7061
rect 570 6810 583 6881
rect 654 6810 670 6881
rect 570 6603 670 6810
rect 570 6532 583 6603
rect 654 6532 670 6603
rect 570 6352 670 6532
rect 570 6281 583 6352
rect 654 6281 670 6352
rect 570 6030 670 6281
rect 570 5959 579 6030
rect 650 5959 670 6030
rect 570 5689 670 5959
rect 570 5618 586 5689
rect 657 5618 670 5689
rect 570 5306 670 5618
rect 570 5235 581 5306
rect 652 5235 670 5306
rect 570 4944 670 5235
rect 570 4873 581 4944
rect 652 4873 670 4944
rect 570 4601 670 4873
rect 570 4530 588 4601
rect 659 4530 670 4601
rect 570 4183 670 4530
rect 570 4112 577 4183
rect 648 4112 670 4183
rect 570 3768 670 4112
rect 570 3697 581 3768
rect 652 3697 670 3768
rect 570 3398 670 3697
rect 570 3327 585 3398
rect 656 3327 670 3398
rect 570 3060 670 3327
rect 1015 7777 1115 7833
rect 1015 7706 1024 7777
rect 1095 7706 1115 7777
rect 1015 7458 1115 7706
rect 1015 7387 1028 7458
rect 1099 7387 1115 7458
rect 1015 7132 1115 7387
rect 1015 7061 1031 7132
rect 1102 7061 1115 7132
rect 1015 6881 1115 7061
rect 1015 6810 1028 6881
rect 1099 6810 1115 6881
rect 1015 6603 1115 6810
rect 1015 6532 1028 6603
rect 1099 6532 1115 6603
rect 1015 6352 1115 6532
rect 1015 6281 1028 6352
rect 1099 6281 1115 6352
rect 1015 6030 1115 6281
rect 1015 5959 1024 6030
rect 1095 5959 1115 6030
rect 1015 5689 1115 5959
rect 1015 5618 1031 5689
rect 1102 5618 1115 5689
rect 1015 5306 1115 5618
rect 1015 5235 1026 5306
rect 1097 5235 1115 5306
rect 1015 4944 1115 5235
rect 1015 4873 1026 4944
rect 1097 4873 1115 4944
rect 1015 4601 1115 4873
rect 1015 4530 1033 4601
rect 1104 4530 1115 4601
rect 1015 4183 1115 4530
rect 1015 4112 1022 4183
rect 1093 4112 1115 4183
rect 1015 3768 1115 4112
rect 1015 3697 1026 3768
rect 1097 3697 1115 3768
rect 1015 3398 1115 3697
rect 1015 3327 1030 3398
rect 1101 3327 1115 3398
rect 1460 7777 1560 8529
rect 1460 7706 1469 7777
rect 1540 7706 1560 7777
rect 1460 7458 1560 7706
rect 1460 7387 1473 7458
rect 1544 7387 1560 7458
rect 1460 7132 1560 7387
rect 1460 7061 1476 7132
rect 1547 7061 1560 7132
rect 1460 6881 1560 7061
rect 1460 6810 1473 6881
rect 1544 6810 1560 6881
rect 1460 6603 1560 6810
rect 1460 6532 1473 6603
rect 1544 6532 1560 6603
rect 1460 6352 1560 6532
rect 1460 6281 1473 6352
rect 1544 6281 1560 6352
rect 1460 6030 1560 6281
rect 1460 5959 1469 6030
rect 1540 5959 1560 6030
rect 1460 5689 1560 5959
rect 1460 5618 1476 5689
rect 1547 5618 1560 5689
rect 1460 5306 1560 5618
rect 1460 5235 1471 5306
rect 1542 5235 1560 5306
rect 1460 4944 1560 5235
rect 1460 4873 1471 4944
rect 1542 4873 1560 4944
rect 1460 4601 1560 4873
rect 1460 4530 1478 4601
rect 1549 4530 1560 4601
rect 1460 4183 1560 4530
rect 1460 4112 1467 4183
rect 1538 4112 1560 4183
rect 1460 3768 1560 4112
rect 1460 3697 1471 3768
rect 1542 3697 1560 3768
rect 1460 3398 1560 3697
rect 1460 3327 1475 3398
rect 1546 3327 1560 3398
rect 1015 3060 1116 3327
rect 1460 3060 1560 3327
rect 1905 7777 2005 7833
rect 1905 7706 1914 7777
rect 1985 7706 2005 7777
rect 1905 7458 2005 7706
rect 1905 7387 1918 7458
rect 1989 7387 2005 7458
rect 1905 7132 2005 7387
rect 1905 7061 1921 7132
rect 1992 7061 2005 7132
rect 1905 6881 2005 7061
rect 1905 6810 1918 6881
rect 1989 6810 2005 6881
rect 1905 6603 2005 6810
rect 1905 6532 1918 6603
rect 1989 6532 2005 6603
rect 1905 6352 2005 6532
rect 1905 6281 1918 6352
rect 1989 6281 2005 6352
rect 1905 6030 2005 6281
rect 1905 5959 1914 6030
rect 1985 5959 2005 6030
rect 1905 5689 2005 5959
rect 1905 5618 1921 5689
rect 1992 5618 2005 5689
rect 1905 5306 2005 5618
rect 1905 5235 1916 5306
rect 1987 5235 2005 5306
rect 1905 4944 2005 5235
rect 1905 4873 1916 4944
rect 1987 4873 2005 4944
rect 1905 4601 2005 4873
rect 1905 4530 1923 4601
rect 1994 4530 2005 4601
rect 1905 4183 2005 4530
rect 1905 4112 1912 4183
rect 1983 4112 2005 4183
rect 1905 3768 2005 4112
rect 1905 3697 1916 3768
rect 1987 3697 2005 3768
rect 1905 3398 2005 3697
rect 1905 3327 1920 3398
rect 1991 3327 2005 3398
rect 2350 7777 2450 8530
rect 2350 7706 2359 7777
rect 2430 7706 2450 7777
rect 2350 7458 2450 7706
rect 2350 7387 2363 7458
rect 2434 7387 2450 7458
rect 2350 7132 2450 7387
rect 2350 7061 2366 7132
rect 2437 7061 2450 7132
rect 2350 6881 2450 7061
rect 2350 6810 2363 6881
rect 2434 6810 2450 6881
rect 2350 6603 2450 6810
rect 2350 6532 2363 6603
rect 2434 6532 2450 6603
rect 2350 6352 2450 6532
rect 2350 6281 2363 6352
rect 2434 6281 2450 6352
rect 2350 6030 2450 6281
rect 2350 5959 2359 6030
rect 2430 5959 2450 6030
rect 2350 5689 2450 5959
rect 2350 5618 2366 5689
rect 2437 5618 2450 5689
rect 2350 5306 2450 5618
rect 2350 5235 2361 5306
rect 2432 5235 2450 5306
rect 2350 4944 2450 5235
rect 2350 4873 2361 4944
rect 2432 4873 2450 4944
rect 2350 4601 2450 4873
rect 2350 4530 2368 4601
rect 2439 4530 2450 4601
rect 2350 4183 2450 4530
rect 2350 4112 2357 4183
rect 2428 4112 2450 4183
rect 2350 3768 2450 4112
rect 2350 3697 2361 3768
rect 2432 3697 2450 3768
rect 2350 3398 2450 3697
rect 2350 3327 2365 3398
rect 2436 3327 2450 3398
rect 1905 3060 2007 3327
rect 2350 3060 2450 3327
rect 2795 7777 2895 7833
rect 2795 7706 2804 7777
rect 2875 7706 2895 7777
rect 2795 7458 2895 7706
rect 2795 7387 2808 7458
rect 2879 7387 2895 7458
rect 2795 7132 2895 7387
rect 2795 7061 2811 7132
rect 2882 7061 2895 7132
rect 2795 6881 2895 7061
rect 2795 6810 2808 6881
rect 2879 6810 2895 6881
rect 2795 6603 2895 6810
rect 2795 6532 2808 6603
rect 2879 6532 2895 6603
rect 2795 6352 2895 6532
rect 2795 6281 2808 6352
rect 2879 6281 2895 6352
rect 2795 6030 2895 6281
rect 2795 5959 2804 6030
rect 2875 5959 2895 6030
rect 2795 5689 2895 5959
rect 2795 5618 2811 5689
rect 2882 5618 2895 5689
rect 2795 5306 2895 5618
rect 2795 5235 2806 5306
rect 2877 5235 2895 5306
rect 2795 4944 2895 5235
rect 2795 4873 2806 4944
rect 2877 4873 2895 4944
rect 2795 4601 2895 4873
rect 2795 4530 2813 4601
rect 2884 4530 2895 4601
rect 2795 4183 2895 4530
rect 2795 4112 2802 4183
rect 2873 4112 2895 4183
rect 2795 3768 2895 4112
rect 2795 3697 2806 3768
rect 2877 3697 2895 3768
rect 2795 3398 2895 3697
rect 2795 3327 2810 3398
rect 2881 3327 2895 3398
rect 2795 3060 2898 3327
rect 640 2521 772 2524
rect 1016 2521 1116 3060
rect 1907 2521 2007 3060
rect 2798 2521 2898 3060
rect -2131 2421 -2111 2521
rect -1637 2421 2898 2521
rect -2131 2406 -2112 2421
rect -2473 2396 -2112 2406
rect -2352 1584 -2252 2396
rect 640 2322 772 2421
rect 640 2279 773 2322
rect 641 2079 773 2279
rect 640 2077 773 2079
rect 640 2000 772 2077
rect 498 1600 898 2000
rect -1003 1185 -603 1193
rect -1003 813 -986 1185
rect -625 813 -603 1185
rect 642 1183 774 1600
rect -248 1083 1654 1183
rect -1003 793 -603 813
rect -237 709 -128 1083
rect -239 606 -127 709
rect 656 696 769 1083
rect 1551 1018 1654 1083
rect 1551 696 1656 1018
rect 224 606 329 664
rect 655 608 769 696
rect 1126 640 1231 643
rect -239 506 -232 606
rect -132 506 -127 606
rect -239 373 -127 506
rect -239 273 -234 373
rect -134 273 -127 373
rect 220 506 228 606
rect 328 506 332 606
rect 220 373 332 506
rect 220 273 226 373
rect 326 273 332 373
rect 655 508 668 608
rect 768 508 769 608
rect 1121 608 1235 640
rect 1121 603 1132 608
rect 655 375 769 508
rect 655 275 666 375
rect 766 275 769 375
rect -239 199 -130 273
rect 220 158 332 273
rect 656 171 769 275
rect 1122 508 1132 603
rect 1232 603 1235 608
rect 1549 610 1661 696
rect 1949 610 2054 643
rect 1232 508 1234 603
rect 1122 375 1234 508
rect 1122 275 1130 375
rect 1230 275 1234 375
rect 1549 510 1558 610
rect 1658 510 1661 610
rect 1549 377 1661 510
rect 1549 277 1556 377
rect 1656 277 1661 377
rect 1944 510 1953 610
rect 2053 510 2056 610
rect 1944 377 2056 510
rect 1944 277 1951 377
rect 2051 277 2056 377
rect 1122 174 1234 275
rect 1551 183 1656 277
rect 224 -171 329 158
rect 1126 -166 1231 174
rect 1944 166 2056 277
rect 1126 -171 1131 -166
rect 224 -174 1131 -171
rect 224 -274 232 -174
rect 332 -266 1131 -174
rect 1949 -166 2054 166
rect 1949 -171 1959 -166
rect 1231 -266 1959 -171
rect 332 -274 2055 -266
rect 224 -276 2055 -274
rect 224 -279 329 -276
<< viali >>
rect -7194 8541 -7024 8711
rect -6351 8538 -6181 8708
rect -5473 8544 -5303 8714
rect -4578 8538 -4408 8708
rect -3729 8547 -3559 8717
rect -1198 8535 -1028 8705
rect -358 8536 -188 8706
rect 538 8546 708 8716
rect 1418 8540 1588 8710
rect 2269 8543 2439 8713
rect 232 -274 332 -174
rect 1131 -266 1231 -166
rect 1959 -266 2059 -166
<< metal1 >>
rect -7397 8717 2743 8985
rect -7397 8714 -3729 8717
rect -7397 8711 -5473 8714
rect -7397 8541 -7194 8711
rect -7024 8708 -5473 8711
rect -7024 8541 -6351 8708
rect -7397 8538 -6351 8541
rect -6181 8544 -5473 8708
rect -5303 8708 -3729 8714
rect -5303 8544 -4578 8708
rect -6181 8538 -4578 8544
rect -4408 8547 -3729 8708
rect -3559 8716 2743 8717
rect -3559 8706 538 8716
rect -3559 8705 -358 8706
rect -3559 8547 -1198 8705
rect -4408 8538 -1198 8547
rect -7397 8535 -1198 8538
rect -1028 8536 -358 8705
rect -188 8546 538 8706
rect 708 8713 2743 8716
rect 708 8710 2269 8713
rect 708 8546 1418 8710
rect -188 8540 1418 8546
rect 1588 8543 2269 8710
rect 2439 8543 2743 8713
rect 1588 8540 2743 8543
rect -188 8536 2743 8540
rect -1028 8535 2743 8536
rect -7397 8393 2743 8535
rect -2301 -166 2153 -98
rect -2301 -174 1131 -166
rect -2301 -274 232 -174
rect 332 -266 1131 -174
rect 1231 -266 1959 -166
rect 2059 -266 2153 -166
rect 332 -274 2153 -266
rect -2301 -355 2153 -274
<< labels >>
flabel metal1 -1033 -239 -1033 -239 0 FreeSans 4000 0 0 0 GND
flabel polycont -807 993 -807 993 0 FreeSans 4000 0 0 0 IN
flabel locali 703 1803 703 1803 0 FreeSans 4000 0 0 0 OUT
flabel metal1 -2357 8674 -2357 8674 0 FreeSans 4000 0 0 0 VDD
flabel locali -2314 1651 -2314 1651 0 FreeSans 4000 0 0 0 A
<< end >>
